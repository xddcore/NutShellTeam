module SRAMTemplate(
  input         clock,
  input         reset,
  output        io_rreq_ready,
  input         io_rreq_valid,
  input  [8:0]  io_rreq_bits_setIdx,
  output [27:0] io_rresp_data_0_tag,
  output [1:0]  io_rresp_data_0__type,
  output [38:0] io_rresp_data_0_target,
  output [2:0]  io_rresp_data_0_brIdx,
  output        io_rresp_data_0_valid,
  input         io_wreq_valid,
  input  [8:0]  io_wreq_bits_setIdx,
  input  [27:0] io_wreq_bits_data_tag,
  input  [1:0]  io_wreq_bits_data__type,
  input  [38:0] io_wreq_bits_data_target,
  input  [2:0]  io_wreq_bits_data_brIdx
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [95:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire [8:0] array_RW0_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_en; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_clk; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmode; // @[SRAMTemplate.scala 76:26]
  wire [72:0] array_RW0_wdata_0; // @[SRAMTemplate.scala 76:26]
  wire [72:0] array_RW0_rdata_0; // @[SRAMTemplate.scala 76:26]
  reg  resetState; // @[SRAMTemplate.scala 80:30]
  reg [8:0] resetSet; // @[Counter.scala 29:33]
  wire  _T_3 = resetSet == 9'h1ff; // @[Counter.scala 38:24]
  wire [8:0] _T_5 = resetSet + 9'h1; // @[Counter.scala 39:22]
  wire  _GEN_1 = resetState & _T_3; // @[Counter.scala 67:17]
  wire  _GEN_2 = _GEN_1 ? 1'h0 : resetState; // @[SRAMTemplate.scala 82:24]
  wire  wen = io_wreq_valid | resetState; // @[SRAMTemplate.scala 88:52]
  wire  _T_6 = ~wen; // @[SRAMTemplate.scala 89:41]
  wire  realRen = io_rreq_valid & _T_6; // @[SRAMTemplate.scala 89:38]
  wire [8:0] setIdx = resetState ? resetSet : io_wreq_bits_setIdx; // @[SRAMTemplate.scala 91:19]
  wire [72:0] _T_11 = {io_wreq_bits_data_tag,io_wreq_bits_data__type,io_wreq_bits_data_target,io_wreq_bits_data_brIdx,1'h1}; // @[SRAMTemplate.scala 92:78]
  reg  _T_20; // @[Hold.scala 28:106]
  reg [72:0] _T_22_0; // @[Reg.scala 27:20]
  wire [72:0] _GEN_14 = _T_20 ? array_RW0_rdata_0 : _T_22_0; // @[Reg.scala 28:19]
  wire  _T_31 = ~resetState; // @[SRAMTemplate.scala 101:21]
  array array ( // @[SRAMTemplate.scala 76:26]
    .RW0_addr(array_RW0_addr),
    .RW0_en(array_RW0_en),
    .RW0_clk(array_RW0_clk),
    .RW0_wmode(array_RW0_wmode),
    .RW0_wdata_0(array_RW0_wdata_0),
    .RW0_rdata_0(array_RW0_rdata_0)
  );
  assign io_rreq_ready = _T_31 & _T_6; // @[SRAMTemplate.scala 101:18]
  assign io_rresp_data_0_tag = _GEN_14[72:45]; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_0__type = _GEN_14[44:43]; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_0_target = _GEN_14[42:4]; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_0_brIdx = _GEN_14[3:1]; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_0_valid = _GEN_14[0]; // @[SRAMTemplate.scala 99:18]
  assign array_RW0_wdata_0 = resetState ? 73'h0 : _T_11;
  assign array_RW0_wmode = io_wreq_valid | resetState;
  assign array_RW0_clk = clock;
  assign array_RW0_en = realRen | wen;
  assign array_RW0_addr = wen ? setIdx : io_rreq_bits_setIdx;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  resetState = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  resetSet = _RAND_1[8:0];
  _RAND_2 = {1{`RANDOM}};
  _T_20 = _RAND_2[0:0];
  _RAND_3 = {3{`RANDOM}};
  _T_22_0 = _RAND_3[72:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    resetState <= reset | _GEN_2;
    if (reset) begin
      resetSet <= 9'h0;
    end else if (resetState) begin
      resetSet <= _T_5;
    end
    _T_20 <= io_rreq_valid & _T_6;
    if (reset) begin
      _T_22_0 <= 73'h0;
    end else if (_T_20) begin
      _T_22_0 <= array_RW0_rdata_0;
    end
  end
endmodule
module BPU_inorder(
  input         clock,
  input         reset,
  input         io_in_pc_valid,
  input  [38:0] io_in_pc_bits,
  output [38:0] io_out_target,
  output        io_out_valid,
  input         io_flush,
  output [2:0]  io_brIdx,
  output        io_crosslineJump,
  input         MOUFlushICache,
  input         bpuUpdateReq_valid,
  input  [38:0] bpuUpdateReq_pc,
  input         bpuUpdateReq_isMissPredict,
  input  [38:0] bpuUpdateReq_actualTarget,
  input         bpuUpdateReq_actualTaken,
  input  [6:0]  bpuUpdateReq_fuOpType,
  input  [1:0]  bpuUpdateReq_btbType,
  input         bpuUpdateReq_isRVC,
  input         MOUFlushTLB
);
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  btb_clock; // @[BPU.scala 302:19]
  wire  btb_reset; // @[BPU.scala 302:19]
  wire  btb_io_rreq_ready; // @[BPU.scala 302:19]
  wire  btb_io_rreq_valid; // @[BPU.scala 302:19]
  wire [8:0] btb_io_rreq_bits_setIdx; // @[BPU.scala 302:19]
  wire [27:0] btb_io_rresp_data_0_tag; // @[BPU.scala 302:19]
  wire [1:0] btb_io_rresp_data_0__type; // @[BPU.scala 302:19]
  wire [38:0] btb_io_rresp_data_0_target; // @[BPU.scala 302:19]
  wire [2:0] btb_io_rresp_data_0_brIdx; // @[BPU.scala 302:19]
  wire  btb_io_rresp_data_0_valid; // @[BPU.scala 302:19]
  wire  btb_io_wreq_valid; // @[BPU.scala 302:19]
  wire [8:0] btb_io_wreq_bits_setIdx; // @[BPU.scala 302:19]
  wire [27:0] btb_io_wreq_bits_data_tag; // @[BPU.scala 302:19]
  wire [1:0] btb_io_wreq_bits_data__type; // @[BPU.scala 302:19]
  wire [38:0] btb_io_wreq_bits_data_target; // @[BPU.scala 302:19]
  wire [2:0] btb_io_wreq_bits_data_brIdx; // @[BPU.scala 302:19]
  reg [1:0] pht [0:511]; // @[BPU.scala 336:16]
  wire [1:0] pht__T_81_data; // @[BPU.scala 336:16]
  wire [8:0] pht__T_81_addr; // @[BPU.scala 336:16]
  wire [1:0] pht__T_139_data; // @[BPU.scala 336:16]
  wire [8:0] pht__T_139_addr; // @[BPU.scala 336:16]
  wire [1:0] pht__T_160_data; // @[BPU.scala 336:16]
  wire [8:0] pht__T_160_addr; // @[BPU.scala 336:16]
  wire  pht__T_160_mask; // @[BPU.scala 336:16]
  wire  pht__T_160_en; // @[BPU.scala 336:16]
  reg [38:0] ras [0:15]; // @[BPU.scala 342:16]
  wire [38:0] ras__T_83_data; // @[BPU.scala 342:16]
  wire [3:0] ras__T_83_addr; // @[BPU.scala 342:16]
  wire [38:0] ras__T_169_data; // @[BPU.scala 342:16]
  wire [3:0] ras__T_169_addr; // @[BPU.scala 342:16]
  wire  ras__T_169_mask; // @[BPU.scala 342:16]
  wire  ras__T_169_en; // @[BPU.scala 342:16]
  reg  flush; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = io_in_pc_valid ? 1'h0 : flush; // @[StopWatch.scala 26:19]
  wire  _GEN_1 = io_flush | _GEN_0; // @[StopWatch.scala 27:20]
  wire  _T_1 = MOUFlushICache | MOUFlushTLB; // @[BPU.scala 308:42]
  reg [38:0] pcLatch; // @[Reg.scala 15:16]
  wire [27:0] btbRead_tag = btb_io_rresp_data_0_tag; // @[BPU.scala 315:21 BPU.scala 316:11]
  wire  _T_27 = btbRead_tag == pcLatch[38:11]; // @[BPU.scala 320:45]
  wire  btbRead_valid = btb_io_rresp_data_0_valid; // @[BPU.scala 315:21 BPU.scala 316:11]
  wire  _T_28 = btbRead_valid & _T_27; // @[BPU.scala 320:30]
  wire  _T_29 = ~flush; // @[BPU.scala 320:76]
  wire  _T_30 = _T_28 & _T_29; // @[BPU.scala 320:73]
  wire  _T_31 = btb_io_rreq_ready & btb_io_rreq_valid; // @[Decoupled.scala 40:37]
  reg  _T_32; // @[BPU.scala 320:93]
  wire  _T_33 = _T_30 & _T_32; // @[BPU.scala 320:83]
  wire [2:0] btbRead_brIdx = btb_io_rresp_data_0_brIdx; // @[BPU.scala 315:21 BPU.scala 316:11]
  wire  _T_36 = pcLatch[1] & btbRead_brIdx[0]; // @[BPU.scala 320:147]
  wire  _T_37 = ~_T_36; // @[BPU.scala 320:134]
  wire  btbHit = _T_33 & _T_37; // @[BPU.scala 320:131]
  wire  crosslineJump = btbRead_brIdx[2] & btbHit; // @[BPU.scala 327:40]
  wire [1:0] _T_64 = io_out_valid ? 2'h3 : 2'h0; // @[Bitwise.scala 72:12]
  reg  phtTaken; // @[Reg.scala 15:16]
  reg [3:0] value; // @[Counter.scala 29:33]
  reg [38:0] rasTarget; // @[Reg.scala 15:16]
  wire  _T_100 = ~bpuUpdateReq_pc[1]; // @[BPU.scala 353:150]
  wire  _T_118 = bpuUpdateReq_pc[2:0] == 3'h6; // @[BPU.scala 367:36]
  wire  _T_119 = ~bpuUpdateReq_isRVC; // @[BPU.scala 367:49]
  wire  _T_120 = _T_118 & _T_119; // @[BPU.scala 367:46]
  wire [1:0] _T_124 = {_T_120,bpuUpdateReq_pc[1]}; // @[Cat.scala 29:58]
  reg [1:0] cnt; // @[BPU.scala 389:20]
  reg  reqLatch_valid; // @[BPU.scala 390:25]
  reg [38:0] reqLatch_pc; // @[BPU.scala 390:25]
  reg  reqLatch_actualTaken; // @[BPU.scala 390:25]
  reg [6:0] reqLatch_fuOpType; // @[BPU.scala 390:25]
  wire  _T_141 = ~reqLatch_fuOpType[3]; // @[ALU.scala 62:30]
  wire  _T_142 = reqLatch_valid & _T_141; // @[BPU.scala 391:24]
  wire [1:0] _T_144 = cnt + 2'h1; // @[BPU.scala 393:33]
  wire [1:0] _T_146 = cnt - 2'h1; // @[BPU.scala 393:44]
  wire  _T_148 = cnt != 2'h3; // @[BPU.scala 394:30]
  wire  _T_149 = reqLatch_actualTaken & _T_148; // @[BPU.scala 394:22]
  wire  _T_150 = ~reqLatch_actualTaken; // @[BPU.scala 394:48]
  wire  _T_151 = cnt != 2'h0; // @[BPU.scala 394:63]
  wire  _T_152 = _T_150 & _T_151; // @[BPU.scala 394:55]
  wire  _T_153 = _T_149 | _T_152; // @[BPU.scala 394:44]
  wire  _T_161 = bpuUpdateReq_fuOpType == 7'h5c; // @[BPU.scala 403:24]
  wire [3:0] _T_163 = value + 4'h1; // @[BPU.scala 404:26]
  wire [38:0] _T_165 = bpuUpdateReq_pc + 39'h2; // @[BPU.scala 404:55]
  wire [38:0] _T_167 = bpuUpdateReq_pc + 39'h4; // @[BPU.scala 404:69]
  wire  _T_172 = bpuUpdateReq_fuOpType == 7'h5e; // @[BPU.scala 408:29]
  wire  _T_173 = value == 4'h0; // @[BPU.scala 409:21]
  wire [3:0] _T_176 = value - 4'h1; // @[BPU.scala 412:53]
  wire [1:0] btbRead__type = btb_io_rresp_data_0__type; // @[BPU.scala 315:21 BPU.scala 316:11]
  wire  _T_178 = btbRead__type == 2'h3; // @[BPU.scala 416:38]
  wire [38:0] btbRead_target = btb_io_rresp_data_0_target; // @[BPU.scala 315:21 BPU.scala 316:11]
  wire [3:0] _T_183 = {1'h1,crosslineJump,_T_64}; // @[Cat.scala 29:58]
  wire [3:0] _GEN_28 = {{1'd0}, btbRead_brIdx}; // @[BPU.scala 419:30]
  wire [3:0] _T_184 = _GEN_28 & _T_183; // @[BPU.scala 419:30]
  wire  _T_185 = btbRead__type == 2'h0; // @[BPU.scala 420:47]
  wire  _T_186 = rasTarget != 39'h0; // @[BPU.scala 420:91]
  wire  _T_188 = _T_185 ? phtTaken : _T_186; // @[BPU.scala 420:32]
  SRAMTemplate btb ( // @[BPU.scala 302:19]
    .clock(btb_clock),
    .reset(btb_reset),
    .io_rreq_ready(btb_io_rreq_ready),
    .io_rreq_valid(btb_io_rreq_valid),
    .io_rreq_bits_setIdx(btb_io_rreq_bits_setIdx),
    .io_rresp_data_0_tag(btb_io_rresp_data_0_tag),
    .io_rresp_data_0__type(btb_io_rresp_data_0__type),
    .io_rresp_data_0_target(btb_io_rresp_data_0_target),
    .io_rresp_data_0_brIdx(btb_io_rresp_data_0_brIdx),
    .io_rresp_data_0_valid(btb_io_rresp_data_0_valid),
    .io_wreq_valid(btb_io_wreq_valid),
    .io_wreq_bits_setIdx(btb_io_wreq_bits_setIdx),
    .io_wreq_bits_data_tag(btb_io_wreq_bits_data_tag),
    .io_wreq_bits_data__type(btb_io_wreq_bits_data__type),
    .io_wreq_bits_data_target(btb_io_wreq_bits_data_target),
    .io_wreq_bits_data_brIdx(btb_io_wreq_bits_data_brIdx)
  );
  assign pht__T_81_addr = io_in_pc_bits[10:2];
  assign pht__T_81_data = pht[pht__T_81_addr]; // @[BPU.scala 336:16]
  assign pht__T_139_addr = bpuUpdateReq_pc[10:2];
  assign pht__T_139_data = pht[pht__T_139_addr]; // @[BPU.scala 336:16]
  assign pht__T_160_data = reqLatch_actualTaken ? _T_144 : _T_146;
  assign pht__T_160_addr = reqLatch_pc[10:2];
  assign pht__T_160_mask = 1'h1;
  assign pht__T_160_en = _T_142 & _T_153;
  assign ras__T_83_addr = value;
  assign ras__T_83_data = ras[ras__T_83_addr]; // @[BPU.scala 342:16]
  assign ras__T_169_data = bpuUpdateReq_isRVC ? _T_165 : _T_167;
  assign ras__T_169_addr = value + 4'h1;
  assign ras__T_169_mask = 1'h1;
  assign ras__T_169_en = bpuUpdateReq_valid & _T_161;
  assign io_out_target = _T_178 ? rasTarget : btbRead_target; // @[BPU.scala 416:17]
  assign io_out_valid = btbHit & _T_188; // @[BPU.scala 420:16]
  assign io_brIdx = _T_184[2:0]; // @[BPU.scala 419:13]
  assign io_crosslineJump = btbRead_brIdx[2] & btbHit; // @[BPU.scala 328:20]
  assign btb_clock = clock;
  assign btb_reset = reset | _T_1; // @[BPU.scala 308:13]
  assign btb_io_rreq_valid = io_in_pc_valid; // @[BPU.scala 311:22]
  assign btb_io_rreq_bits_setIdx = io_in_pc_bits[10:2]; // @[BPU.scala 312:28]
  assign btb_io_wreq_valid = bpuUpdateReq_isMissPredict & bpuUpdateReq_valid; // @[BPU.scala 375:22]
  assign btb_io_wreq_bits_setIdx = bpuUpdateReq_pc[10:2]; // @[BPU.scala 376:28]
  assign btb_io_wreq_bits_data_tag = bpuUpdateReq_pc[38:11]; // @[BPU.scala 377:26]
  assign btb_io_wreq_bits_data__type = bpuUpdateReq_btbType; // @[BPU.scala 377:26]
  assign btb_io_wreq_bits_data_target = bpuUpdateReq_actualTarget; // @[BPU.scala 377:26]
  assign btb_io_wreq_bits_data_brIdx = {_T_124,_T_100}; // @[BPU.scala 377:26]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 512; initvar = initvar+1)
    pht[initvar] = _RAND_0[1:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    ras[initvar] = _RAND_1[38:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  flush = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  pcLatch = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  _T_32 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  phtTaken = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  value = _RAND_6[3:0];
  _RAND_7 = {2{`RANDOM}};
  rasTarget = _RAND_7[38:0];
  _RAND_8 = {1{`RANDOM}};
  cnt = _RAND_8[1:0];
  _RAND_9 = {1{`RANDOM}};
  reqLatch_valid = _RAND_9[0:0];
  _RAND_10 = {2{`RANDOM}};
  reqLatch_pc = _RAND_10[38:0];
  _RAND_11 = {1{`RANDOM}};
  reqLatch_actualTaken = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  reqLatch_fuOpType = _RAND_12[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(pht__T_160_en & pht__T_160_mask) begin
      pht[pht__T_160_addr] <= pht__T_160_data; // @[BPU.scala 336:16]
    end
    if(ras__T_169_en & ras__T_169_mask) begin
      ras[ras__T_169_addr] <= ras__T_169_data; // @[BPU.scala 342:16]
    end
    if (reset) begin
      flush <= 1'h0;
    end else begin
      flush <= _GEN_1;
    end
    if (io_in_pc_valid) begin
      pcLatch <= io_in_pc_bits;
    end
    if (reset) begin
      _T_32 <= 1'h0;
    end else begin
      _T_32 <= _T_31;
    end
    if (io_in_pc_valid) begin
      phtTaken <= pht__T_81_data[1];
    end
    if (reset) begin
      value <= 4'h0;
    end else if (bpuUpdateReq_valid) begin
      if (_T_161) begin
        value <= _T_163;
      end else if (_T_172) begin
        if (_T_173) begin
          value <= 4'h0;
        end else begin
          value <= _T_176;
        end
      end
    end
    if (io_in_pc_valid) begin
      rasTarget <= ras__T_83_data;
    end
    cnt <= pht__T_139_data;
    reqLatch_valid <= bpuUpdateReq_valid;
    reqLatch_pc <= bpuUpdateReq_pc;
    reqLatch_actualTaken <= bpuUpdateReq_actualTaken;
    reqLatch_fuOpType <= bpuUpdateReq_fuOpType;
  end
endmodule
module IFU_inorder(
  input         clock,
  input         reset,
  input         io_imem_req_ready,
  output        io_imem_req_valid,
  output [38:0] io_imem_req_bits_addr,
  output [81:0] io_imem_req_bits_user,
  output        io_imem_resp_ready,
  input         io_imem_resp_valid,
  input  [63:0] io_imem_resp_bits_rdata,
  input  [81:0] io_imem_resp_bits_user,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_instr,
  output [38:0] io_out_bits_pc,
  output [38:0] io_out_bits_pnpc,
  output        io_out_bits_exceptionVec_12,
  output [3:0]  io_out_bits_brIdx,
  input  [38:0] io_redirect_target,
  input         io_redirect_valid,
  output [3:0]  io_flushVec,
  input         io_ipf,
  input         flushICache,
  input         _T_243_valid,
  input  [38:0] _T_243_pc,
  input         _T_243_isMissPredict,
  input  [38:0] _T_243_actualTarget,
  input         _T_243_actualTaken,
  input  [6:0]  _T_243_fuOpType,
  input  [1:0]  _T_243_btbType,
  input         _T_243_isRVC,
  input         flushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  wire  bp1_clock; // @[IFU.scala 325:19]
  wire  bp1_reset; // @[IFU.scala 325:19]
  wire  bp1_io_in_pc_valid; // @[IFU.scala 325:19]
  wire [38:0] bp1_io_in_pc_bits; // @[IFU.scala 325:19]
  wire [38:0] bp1_io_out_target; // @[IFU.scala 325:19]
  wire  bp1_io_out_valid; // @[IFU.scala 325:19]
  wire  bp1_io_flush; // @[IFU.scala 325:19]
  wire [2:0] bp1_io_brIdx; // @[IFU.scala 325:19]
  wire  bp1_io_crosslineJump; // @[IFU.scala 325:19]
  wire  bp1_MOUFlushICache; // @[IFU.scala 325:19]
  wire  bp1_bpuUpdateReq_valid; // @[IFU.scala 325:19]
  wire [38:0] bp1_bpuUpdateReq_pc; // @[IFU.scala 325:19]
  wire  bp1_bpuUpdateReq_isMissPredict; // @[IFU.scala 325:19]
  wire [38:0] bp1_bpuUpdateReq_actualTarget; // @[IFU.scala 325:19]
  wire  bp1_bpuUpdateReq_actualTaken; // @[IFU.scala 325:19]
  wire [6:0] bp1_bpuUpdateReq_fuOpType; // @[IFU.scala 325:19]
  wire [1:0] bp1_bpuUpdateReq_btbType; // @[IFU.scala 325:19]
  wire  bp1_bpuUpdateReq_isRVC; // @[IFU.scala 325:19]
  wire  bp1_MOUFlushTLB; // @[IFU.scala 325:19]
  reg [38:0] pc; // @[IFU.scala 321:19]
  wire  _T = io_imem_req_ready & io_imem_req_valid; // @[Decoupled.scala 40:37]
  wire  pcUpdate = io_redirect_valid | _T; // @[IFU.scala 322:36]
  wire [38:0] _T_3 = pc + 39'h2; // @[IFU.scala 323:28]
  wire [38:0] _T_5 = pc + 39'h4; // @[IFU.scala 323:38]
  wire [38:0] snpc = pc[1] ? _T_3 : _T_5; // @[IFU.scala 323:17]
  reg  crosslineJumpLatch; // @[IFU.scala 328:35]
  wire  _T_6 = pcUpdate | bp1_io_flush; // @[IFU.scala 329:17]
  wire  _T_7 = ~crosslineJumpLatch; // @[IFU.scala 330:71]
  wire  _T_8 = bp1_io_crosslineJump & _T_7; // @[IFU.scala 330:68]
  reg [38:0] crosslineJumpTarget; // @[Reg.scala 15:16]
  wire [38:0] pnpc = bp1_io_crosslineJump ? snpc : bp1_io_out_target; // @[IFU.scala 337:17]
  wire [38:0] _T_11 = bp1_io_out_valid ? pnpc : snpc; // @[IFU.scala 339:104]
  wire [38:0] _T_12 = crosslineJumpLatch ? crosslineJumpTarget : _T_11; // @[IFU.scala 339:59]
  wire [38:0] npc = io_redirect_valid ? io_redirect_target : _T_12; // @[IFU.scala 339:16]
  wire  _T_13 = bp1_io_out_valid ? 1'h0 : 1'h1; // @[IFU.scala 340:114]
  wire  _T_14 = bp1_io_crosslineJump | _T_13; // @[IFU.scala 340:87]
  wire  _T_15 = crosslineJumpLatch ? 1'h0 : _T_14; // @[IFU.scala 340:54]
  wire  npcIsSeq = io_redirect_valid ? 1'h0 : _T_15; // @[IFU.scala 340:21]
  wire [2:0] _T_16 = io_redirect_valid ? 3'h0 : bp1_io_brIdx; // @[IFU.scala 348:29]
  wire [42:0] _T_34 = {npcIsSeq,_T_16,npc}; // @[Cat.scala 29:58]
  wire  _T_62 = ~io_flushVec[0]; // @[IFU.scala 390:41]
  wire  _T_64 = io_imem_resp_ready & io_imem_resp_valid; // @[Decoupled.scala 40:37]
  reg  _T_65; // @[StopWatch.scala 24:20]
  wire  _GEN_3 = io_imem_req_valid | _T_65; // @[StopWatch.scala 30:20]
  wire  _T_66 = |io_flushVec; // @[IFU.scala 393:37]
  BPU_inorder bp1 ( // @[IFU.scala 325:19]
    .clock(bp1_clock),
    .reset(bp1_reset),
    .io_in_pc_valid(bp1_io_in_pc_valid),
    .io_in_pc_bits(bp1_io_in_pc_bits),
    .io_out_target(bp1_io_out_target),
    .io_out_valid(bp1_io_out_valid),
    .io_flush(bp1_io_flush),
    .io_brIdx(bp1_io_brIdx),
    .io_crosslineJump(bp1_io_crosslineJump),
    .MOUFlushICache(bp1_MOUFlushICache),
    .bpuUpdateReq_valid(bp1_bpuUpdateReq_valid),
    .bpuUpdateReq_pc(bp1_bpuUpdateReq_pc),
    .bpuUpdateReq_isMissPredict(bp1_bpuUpdateReq_isMissPredict),
    .bpuUpdateReq_actualTarget(bp1_bpuUpdateReq_actualTarget),
    .bpuUpdateReq_actualTaken(bp1_bpuUpdateReq_actualTaken),
    .bpuUpdateReq_fuOpType(bp1_bpuUpdateReq_fuOpType),
    .bpuUpdateReq_btbType(bp1_bpuUpdateReq_btbType),
    .bpuUpdateReq_isRVC(bp1_bpuUpdateReq_isRVC),
    .MOUFlushTLB(bp1_MOUFlushTLB)
  );
  assign io_imem_req_valid = io_out_ready; // @[IFU.scala 371:21]
  assign io_imem_req_bits_addr = {pc[38:1],1'h0}; // @[SimpleBus.scala 64:15]
  assign io_imem_req_bits_user = {_T_34,pc}; // @[SimpleBus.scala 69:21]
  assign io_imem_resp_ready = io_out_ready | io_flushVec[0]; // @[IFU.scala 373:22]
  assign io_out_valid = io_imem_resp_valid & _T_62; // @[IFU.scala 390:16]
  assign io_out_bits_instr = io_imem_resp_bits_rdata; // @[IFU.scala 383:21]
  assign io_out_bits_pc = io_imem_resp_bits_user[38:0]; // @[IFU.scala 385:20]
  assign io_out_bits_pnpc = io_imem_resp_bits_user[77:39]; // @[IFU.scala 386:22]
  assign io_out_bits_exceptionVec_12 = io_ipf; // @[IFU.scala 389:44]
  assign io_out_bits_brIdx = io_imem_resp_bits_user[81:78]; // @[IFU.scala 387:23]
  assign io_flushVec = io_redirect_valid ? 4'hf : 4'h0; // @[IFU.scala 366:15]
  assign bp1_clock = clock;
  assign bp1_reset = reset;
  assign bp1_io_in_pc_valid = io_imem_req_ready & io_imem_req_valid; // @[IFU.scala 351:22]
  assign bp1_io_in_pc_bits = io_redirect_valid ? io_redirect_target : _T_12; // @[IFU.scala 352:21]
  assign bp1_io_flush = io_redirect_valid; // @[IFU.scala 357:16]
  assign bp1_MOUFlushICache = flushICache;
  assign bp1_bpuUpdateReq_valid = _T_243_valid;
  assign bp1_bpuUpdateReq_pc = _T_243_pc;
  assign bp1_bpuUpdateReq_isMissPredict = _T_243_isMissPredict;
  assign bp1_bpuUpdateReq_actualTarget = _T_243_actualTarget;
  assign bp1_bpuUpdateReq_actualTaken = _T_243_actualTaken;
  assign bp1_bpuUpdateReq_fuOpType = _T_243_fuOpType;
  assign bp1_bpuUpdateReq_btbType = _T_243_btbType;
  assign bp1_bpuUpdateReq_isRVC = _T_243_isRVC;
  assign bp1_MOUFlushTLB = flushTLB;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  pc = _RAND_0[38:0];
  _RAND_1 = {1{`RANDOM}};
  crosslineJumpLatch = _RAND_1[0:0];
  _RAND_2 = {2{`RANDOM}};
  crosslineJumpTarget = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  _T_65 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      pc <= 39'h60000000;
    end else if (pcUpdate) begin
      if (io_redirect_valid) begin
        pc <= io_redirect_target;
      end else if (crosslineJumpLatch) begin
        pc <= crosslineJumpTarget;
      end else if (bp1_io_out_valid) begin
        if (bp1_io_crosslineJump) begin
          if (pc[1]) begin
            pc <= _T_3;
          end else begin
            pc <= _T_5;
          end
        end else begin
          pc <= bp1_io_out_target;
        end
      end else if (pc[1]) begin
        pc <= _T_3;
      end else begin
        pc <= _T_5;
      end
    end
    if (reset) begin
      crosslineJumpLatch <= 1'h0;
    end else if (_T_6) begin
      if (bp1_io_flush) begin
        crosslineJumpLatch <= 1'h0;
      end else begin
        crosslineJumpLatch <= _T_8;
      end
    end
    if (bp1_io_crosslineJump) begin
      crosslineJumpTarget <= bp1_io_out_target;
    end
    if (reset) begin
      _T_65 <= 1'h0;
    end else if (_T_64) begin
      _T_65 <= 1'h0;
    end else begin
      _T_65 <= _GEN_3;
    end
  end
endmodule
module NaiveRVCAlignBuffer(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_instr,
  input  [38:0] io_in_bits_pc,
  input  [38:0] io_in_bits_pnpc,
  input         io_in_bits_exceptionVec_12,
  input  [3:0]  io_in_bits_brIdx,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_instr,
  output [38:0] io_out_bits_pc,
  output [38:0] io_out_bits_pnpc,
  output        io_out_bits_exceptionVec_12,
  output [3:0]  io_out_bits_brIdx,
  output        io_out_bits_crossPageIPFFix,
  input         io_flush
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[NaiveIBF.scala 39:22]
  wire  _T_83 = state == 2'h2; // @[NaiveIBF.scala 90:23]
  wire  _T_84 = state == 2'h3; // @[NaiveIBF.scala 90:47]
  wire  _T_85 = _T_83 | _T_84; // @[NaiveIBF.scala 90:38]
  wire [79:0] instIn = {16'h0,io_in_bits_instr}; // @[Cat.scala 29:58]
  reg [15:0] specialInstR; // @[NaiveIBF.scala 66:25]
  wire [31:0] _T_87 = {instIn[15:0],specialInstR}; // @[Cat.scala 29:58]
  wire  _T_1 = state == 2'h0; // @[NaiveIBF.scala 41:28]
  reg [2:0] pcOffsetR; // @[NaiveIBF.scala 40:26]
  wire [2:0] pcOffset = _T_1 ? io_in_bits_pc[2:0] : pcOffsetR; // @[NaiveIBF.scala 41:21]
  wire  _T_92 = 3'h0 == pcOffset; // @[LookupTree.scala 24:34]
  wire [31:0] _T_96 = _T_92 ? instIn[31:0] : 32'h0; // @[Mux.scala 27:72]
  wire  _T_93 = 3'h2 == pcOffset; // @[LookupTree.scala 24:34]
  wire [31:0] _T_97 = _T_93 ? instIn[47:16] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_100 = _T_96 | _T_97; // @[Mux.scala 27:72]
  wire  _T_94 = 3'h4 == pcOffset; // @[LookupTree.scala 24:34]
  wire [31:0] _T_98 = _T_94 ? instIn[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_101 = _T_100 | _T_98; // @[Mux.scala 27:72]
  wire  _T_95 = 3'h6 == pcOffset; // @[LookupTree.scala 24:34]
  wire [31:0] _T_99 = _T_95 ? instIn[79:48] : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_102 = _T_101 | _T_99; // @[Mux.scala 27:72]
  wire [31:0] instr = _T_85 ? _T_87 : _T_102; // @[NaiveIBF.scala 90:15]
  wire  isRVC = instr[1:0] != 2'h3; // @[NaiveIBF.scala 34:26]
  wire  _T_3 = pcOffset == 3'h0; // @[NaiveIBF.scala 48:28]
  wire  _T_4 = ~isRVC; // @[NaiveIBF.scala 48:40]
  wire  _T_6 = _T_4 | io_in_bits_brIdx[0]; // @[NaiveIBF.scala 48:47]
  wire  _T_7 = _T_3 & _T_6; // @[NaiveIBF.scala 48:36]
  wire  _T_8 = pcOffset == 3'h4; // @[NaiveIBF.scala 48:72]
  wire  _T_12 = _T_8 & _T_6; // @[NaiveIBF.scala 48:80]
  wire  _T_13 = _T_7 | _T_12; // @[NaiveIBF.scala 48:60]
  wire  _T_14 = pcOffset == 3'h2; // @[NaiveIBF.scala 48:116]
  wire  _T_16 = isRVC | io_in_bits_brIdx[1]; // @[NaiveIBF.scala 48:134]
  wire  _T_17 = _T_14 & _T_16; // @[NaiveIBF.scala 48:124]
  wire  _T_18 = _T_13 | _T_17; // @[NaiveIBF.scala 48:104]
  wire  _T_19 = pcOffset == 3'h6; // @[NaiveIBF.scala 48:159]
  wire  _T_20 = _T_19 & isRVC; // @[NaiveIBF.scala 48:167]
  wire  rvcFinish = _T_18 | _T_20; // @[NaiveIBF.scala 48:147]
  wire  _T_23 = ~io_in_bits_brIdx[0]; // @[NaiveIBF.scala 51:47]
  wire  _T_24 = isRVC & _T_23; // @[NaiveIBF.scala 51:44]
  wire  _T_25 = _T_3 & _T_24; // @[NaiveIBF.scala 51:34]
  wire  _T_30 = _T_8 & _T_24; // @[NaiveIBF.scala 51:78]
  wire  _T_31 = _T_25 | _T_30; // @[NaiveIBF.scala 51:58]
  wire  _T_34 = _T_14 & _T_4; // @[NaiveIBF.scala 51:122]
  wire  _T_36 = ~io_in_bits_brIdx[1]; // @[NaiveIBF.scala 51:135]
  wire  _T_37 = _T_34 & _T_36; // @[NaiveIBF.scala 51:132]
  wire  rvcNext = _T_31 | _T_37; // @[NaiveIBF.scala 51:102]
  wire  _T_40 = _T_19 & _T_4; // @[NaiveIBF.scala 52:37]
  wire  _T_42 = ~io_in_bits_brIdx[2]; // @[NaiveIBF.scala 52:50]
  wire  rvcSpecial = _T_40 & _T_42; // @[NaiveIBF.scala 52:47]
  wire  rvcSpecialJump = _T_40 & io_in_bits_brIdx[2]; // @[NaiveIBF.scala 53:51]
  wire  pnpcIsSeq = io_in_bits_brIdx[3]; // @[NaiveIBF.scala 54:24]
  wire  _T_48 = state == 2'h1; // @[NaiveIBF.scala 57:45]
  wire  _T_49 = _T_1 | _T_48; // @[NaiveIBF.scala 57:36]
  wire  _T_50 = _T_49 & rvcSpecial; // @[NaiveIBF.scala 57:58]
  wire  _T_51 = _T_50 & io_in_valid; // @[NaiveIBF.scala 57:72]
  wire  _T_52 = ~pnpcIsSeq; // @[NaiveIBF.scala 57:90]
  wire  flushIFU = _T_51 & _T_52; // @[NaiveIBF.scala 57:87]
  wire  _T_62 = ~flushIFU; // @[NaiveIBF.scala 59:10]
  wire  _T_64 = _T_62 | reset; // @[NaiveIBF.scala 59:9]
  wire  _T_65 = ~_T_64; // @[NaiveIBF.scala 59:9]
  wire  _T_69 = rvcSpecial | rvcSpecialJump; // @[NaiveIBF.scala 60:81]
  wire  _T_70 = _T_49 & _T_69; // @[NaiveIBF.scala 60:66]
  wire  _T_71 = _T_70 & io_in_valid; // @[NaiveIBF.scala 60:100]
  wire  loadNextInstline = _T_71 & pnpcIsSeq; // @[NaiveIBF.scala 60:115]
  reg [38:0] specialPCR; // @[NaiveIBF.scala 64:23]
  reg [38:0] specialNPCR; // @[NaiveIBF.scala 65:24]
  reg  specialIPFR; // @[NaiveIBF.scala 67:28]
  wire  _T_79 = io_in_bits_pnpc[2:0] == 3'h4; // @[NaiveIBF.scala 69:78]
  wire  _T_80 = _T_34 & _T_79; // @[NaiveIBF.scala 69:54]
  wire  rvcForceLoadNext = _T_80 & _T_36; // @[NaiveIBF.scala 69:86]
  wire  _T_105 = ~io_flush; // @[NaiveIBF.scala 97:8]
  wire  _T_106 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_107 = rvcFinish | rvcNext; // @[NaiveIBF.scala 100:28]
  wire  _T_108 = rvcFinish | rvcForceLoadNext; // @[NaiveIBF.scala 101:28]
  wire [38:0] _T_110 = io_in_bits_pc + 39'h2; // @[NaiveIBF.scala 103:76]
  wire [38:0] _T_112 = io_in_bits_pc + 39'h4; // @[NaiveIBF.scala 103:95]
  wire [38:0] _T_113 = isRVC ? _T_110 : _T_112; // @[NaiveIBF.scala 103:55]
  wire [38:0] _T_114 = rvcFinish ? io_in_bits_pnpc : _T_113; // @[NaiveIBF.scala 103:23]
  wire  _T_115 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_116 = _T_115 & rvcFinish; // @[NaiveIBF.scala 104:28]
  wire  _T_118 = _T_115 & rvcNext; // @[NaiveIBF.scala 105:28]
  wire [2:0] _T_119 = isRVC ? 3'h2 : 3'h4; // @[NaiveIBF.scala 107:38]
  wire [2:0] _T_121 = pcOffset + _T_119; // @[NaiveIBF.scala 107:33]
  wire  _T_122 = rvcSpecial & io_in_valid; // @[NaiveIBF.scala 109:25]
  wire  _T_126 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire [38:0] _T_131 = {io_in_bits_pc[38:3],pcOffsetR}; // @[Cat.scala 29:58]
  wire  _T_149 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_153 = 2'h3 == state; // @[Conditional.scala 37:30]
  wire [38:0] _GEN_27 = _T_153 ? specialPCR : 39'h0; // @[Conditional.scala 39:67]
  wire [38:0] _GEN_32 = _T_149 ? specialPCR : _GEN_27; // @[Conditional.scala 39:67]
  wire [38:0] _GEN_40 = _T_126 ? _T_131 : _GEN_32; // @[Conditional.scala 39:67]
  wire [38:0] pcOut = _T_106 ? io_in_bits_pc : _GEN_40; // @[Conditional.scala 40:58]
  wire  _T_124 = rvcSpecialJump & io_in_valid; // @[NaiveIBF.scala 115:29]
  wire [38:0] _T_133 = pcOut + 39'h2; // @[NaiveIBF.scala 127:68]
  wire [38:0] _T_135 = pcOut + 39'h4; // @[NaiveIBF.scala 127:79]
  wire [38:0] _T_136 = isRVC ? _T_133 : _T_135; // @[NaiveIBF.scala 127:55]
  wire [38:0] _T_137 = rvcFinish ? io_in_bits_pnpc : _T_136; // @[NaiveIBF.scala 127:23]
  wire [38:0] _T_151 = specialPCR + 39'h4; // @[NaiveIBF.scala 150:31]
  wire [38:0] _GEN_28 = _T_153 ? specialNPCR : 39'h0; // @[Conditional.scala 39:67]
  wire  _GEN_29 = _T_153 & io_in_valid; // @[Conditional.scala 39:67]
  wire [38:0] _GEN_33 = _T_149 ? _T_151 : _GEN_28; // @[Conditional.scala 39:67]
  wire  _GEN_34 = _T_149 ? io_in_valid : _GEN_29; // @[Conditional.scala 39:67]
  wire  _GEN_35 = _T_149 ? 1'h0 : _T_153; // @[Conditional.scala 39:67]
  wire  _GEN_38 = _T_126 ? _T_107 : _GEN_34; // @[Conditional.scala 39:67]
  wire  _GEN_39 = _T_126 ? _T_108 : _GEN_35; // @[Conditional.scala 39:67]
  wire [38:0] _GEN_41 = _T_126 ? _T_137 : _GEN_33; // @[Conditional.scala 39:67]
  wire  canGo = _T_106 ? _T_107 : _GEN_38; // @[Conditional.scala 40:58]
  wire  canIn = _T_106 ? _T_108 : _GEN_39; // @[Conditional.scala 40:58]
  wire [38:0] pnpcOut = _T_106 ? _T_114 : _GEN_41; // @[Conditional.scala 40:58]
  wire  _T_157 = pnpcOut == _T_135; // @[NaiveIBF.scala 185:37]
  wire  _T_159 = _T_157 & _T_4; // @[NaiveIBF.scala 185:51]
  wire  _T_162 = pnpcOut == _T_133; // @[NaiveIBF.scala 185:74]
  wire  _T_163 = _T_162 & isRVC; // @[NaiveIBF.scala 185:88]
  wire  _T_164 = _T_159 | _T_163; // @[NaiveIBF.scala 185:62]
  wire  _T_165 = _T_164 ? 1'h0 : 1'h1; // @[NaiveIBF.scala 185:27]
  wire  _T_167 = ~io_in_valid; // @[NaiveIBF.scala 188:19]
  wire  _T_169 = _T_115 & canIn; // @[NaiveIBF.scala 188:50]
  wire  _T_170 = _T_167 | _T_169; // @[NaiveIBF.scala 188:32]
  wire  _T_174 = _T_84 | _T_83; // @[NaiveIBF.scala 191:133]
  wire  _T_175 = specialIPFR & _T_174; // @[NaiveIBF.scala 191:102]
  wire  _T_180 = io_in_bits_exceptionVec_12 & _T_174; // @[NaiveIBF.scala 192:74]
  wire  _T_181 = ~specialIPFR; // @[NaiveIBF.scala 192:133]
  assign io_in_ready = _T_170 | loadNextInstline; // @[NaiveIBF.scala 188:15]
  assign io_out_valid = io_in_valid & canGo; // @[NaiveIBF.scala 187:16]
  assign io_out_bits_instr = {{32'd0}, instr}; // @[NaiveIBF.scala 184:21]
  assign io_out_bits_pc = _T_106 ? io_in_bits_pc : _GEN_40; // @[NaiveIBF.scala 182:18]
  assign io_out_bits_pnpc = _T_106 ? _T_114 : _GEN_41; // @[NaiveIBF.scala 183:20]
  assign io_out_bits_exceptionVec_12 = io_in_bits_exceptionVec_12 | _T_175; // @[NaiveIBF.scala 190:28 NaiveIBF.scala 191:44]
  assign io_out_bits_brIdx = {{3'd0}, _T_165}; // @[NaiveIBF.scala 185:21]
  assign io_out_bits_crossPageIPFFix = _T_180 & _T_181; // @[NaiveIBF.scala 192:31]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  specialInstR = _RAND_1[15:0];
  _RAND_2 = {1{`RANDOM}};
  pcOffsetR = _RAND_2[2:0];
  _RAND_3 = {2{`RANDOM}};
  specialPCR = _RAND_3[38:0];
  _RAND_4 = {2{`RANDOM}};
  specialNPCR = _RAND_4[38:0];
  _RAND_5 = {1{`RANDOM}};
  specialIPFR = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else if (_T_105) begin
      if (_T_106) begin
        if (_T_124) begin
          state <= 2'h3;
        end else if (_T_122) begin
          state <= 2'h2;
        end else if (_T_118) begin
          state <= 2'h1;
        end else if (_T_116) begin
          state <= 2'h0;
        end
      end else if (_T_126) begin
        if (_T_124) begin
          state <= 2'h3;
        end else if (_T_122) begin
          state <= 2'h2;
        end else if (_T_118) begin
          state <= 2'h1;
        end else if (_T_116) begin
          state <= 2'h0;
        end
      end else if (_T_149) begin
        if (_T_115) begin
          state <= 2'h1;
        end
      end else if (_T_153) begin
        if (_T_115) begin
          state <= 2'h0;
        end
      end
    end else begin
      state <= 2'h0;
    end
    if (_T_105) begin
      if (_T_106) begin
        if (_T_124) begin
          specialInstR <= io_in_bits_instr[63:48];
        end else if (_T_122) begin
          specialInstR <= io_in_bits_instr[63:48];
        end
      end else if (_T_126) begin
        if (_T_124) begin
          specialInstR <= io_in_bits_instr[63:48];
        end else if (_T_122) begin
          specialInstR <= io_in_bits_instr[63:48];
        end
      end
    end
    if (reset) begin
      pcOffsetR <= 3'h0;
    end else if (_T_105) begin
      if (_T_106) begin
        if (_T_118) begin
          pcOffsetR <= _T_121;
        end
      end else if (_T_126) begin
        if (_T_118) begin
          pcOffsetR <= _T_121;
        end
      end else if (_T_149) begin
        if (_T_115) begin
          pcOffsetR <= 3'h2;
        end
      end
    end
    if (_T_105) begin
      if (_T_106) begin
        if (_T_124) begin
          if (_T_106) begin
            specialPCR <= io_in_bits_pc;
          end else if (_T_126) begin
            specialPCR <= _T_131;
          end else if (!(_T_149)) begin
            if (!(_T_153)) begin
              specialPCR <= 39'h0;
            end
          end
        end else if (_T_122) begin
          if (_T_106) begin
            specialPCR <= io_in_bits_pc;
          end else if (_T_126) begin
            specialPCR <= _T_131;
          end else if (!(_T_149)) begin
            if (!(_T_153)) begin
              specialPCR <= 39'h0;
            end
          end
        end
      end else if (_T_126) begin
        if (_T_124) begin
          if (_T_106) begin
            specialPCR <= io_in_bits_pc;
          end else if (_T_126) begin
            specialPCR <= _T_131;
          end else if (!(_T_149)) begin
            if (!(_T_153)) begin
              specialPCR <= 39'h0;
            end
          end
        end else if (_T_122) begin
          if (_T_106) begin
            specialPCR <= io_in_bits_pc;
          end else if (_T_126) begin
            specialPCR <= _T_131;
          end else if (!(_T_149)) begin
            if (!(_T_153)) begin
              specialPCR <= 39'h0;
            end
          end
        end
      end
    end
    if (_T_105) begin
      if (_T_106) begin
        if (_T_124) begin
          specialNPCR <= io_in_bits_pnpc;
        end
      end else if (_T_126) begin
        if (_T_124) begin
          specialNPCR <= io_in_bits_pnpc;
        end
      end
    end
    if (reset) begin
      specialIPFR <= 1'h0;
    end else if (_T_105) begin
      if (_T_106) begin
        if (_T_124) begin
          specialIPFR <= io_in_bits_exceptionVec_12;
        end else if (_T_122) begin
          specialIPFR <= io_in_bits_exceptionVec_12;
        end
      end else if (_T_126) begin
        if (_T_124) begin
          specialIPFR <= io_in_bits_exceptionVec_12;
        end else if (_T_122) begin
          specialIPFR <= io_in_bits_exceptionVec_12;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_65) begin
          $fwrite(32'h80000002,"Assertion failed\n    at NaiveIBF.scala:59 assert(!flushIFU)\n"); // @[NaiveIBF.scala 59:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_65) begin
          $fatal; // @[NaiveIBF.scala 59:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Decoder(
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_instr,
  input  [38:0] io_in_bits_pc,
  input  [38:0] io_in_bits_pnpc,
  input         io_in_bits_exceptionVec_12,
  input  [3:0]  io_in_bits_brIdx,
  input         io_in_bits_crossPageIPFFix,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_cf_instr,
  output [38:0] io_out_bits_cf_pc,
  output [38:0] io_out_bits_cf_pnpc,
  output        io_out_bits_cf_exceptionVec_1,
  output        io_out_bits_cf_exceptionVec_2,
  output        io_out_bits_cf_exceptionVec_12,
  output        io_out_bits_cf_intrVec_0,
  output        io_out_bits_cf_intrVec_1,
  output        io_out_bits_cf_intrVec_2,
  output        io_out_bits_cf_intrVec_3,
  output        io_out_bits_cf_intrVec_4,
  output        io_out_bits_cf_intrVec_5,
  output        io_out_bits_cf_intrVec_6,
  output        io_out_bits_cf_intrVec_7,
  output        io_out_bits_cf_intrVec_8,
  output        io_out_bits_cf_intrVec_9,
  output        io_out_bits_cf_intrVec_10,
  output        io_out_bits_cf_intrVec_11,
  output [3:0]  io_out_bits_cf_brIdx,
  output        io_out_bits_cf_crossPageIPFFix,
  output        io_out_bits_ctrl_src1Type,
  output        io_out_bits_ctrl_src2Type,
  output [2:0]  io_out_bits_ctrl_fuType,
  output [6:0]  io_out_bits_ctrl_fuOpType,
  output [4:0]  io_out_bits_ctrl_rfSrc1,
  output [4:0]  io_out_bits_ctrl_rfSrc2,
  output        io_out_bits_ctrl_rfWen,
  output [4:0]  io_out_bits_ctrl_rfDest,
  output [63:0] io_out_bits_data_imm,
  input         DTLBENABLE,
  input  [11:0] intrVecIDU
);
  wire [63:0] _T = io_in_bits_instr & 64'h707f; // @[Lookup.scala 31:38]
  wire  _T_1 = 64'h13 == _T; // @[Lookup.scala 31:38]
  wire [63:0] _T_2 = io_in_bits_instr & 64'hfc00707f; // @[Lookup.scala 31:38]
  wire  _T_3 = 64'h1013 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_5 = 64'h2013 == _T; // @[Lookup.scala 31:38]
  wire  _T_7 = 64'h3013 == _T; // @[Lookup.scala 31:38]
  wire  _T_9 = 64'h4013 == _T; // @[Lookup.scala 31:38]
  wire  _T_11 = 64'h5013 == _T_2; // @[Lookup.scala 31:38]
  wire  _T_13 = 64'h6013 == _T; // @[Lookup.scala 31:38]
  wire  _T_15 = 64'h7013 == _T; // @[Lookup.scala 31:38]
  wire  _T_17 = 64'h40005013 == _T_2; // @[Lookup.scala 31:38]
  wire [63:0] _T_18 = io_in_bits_instr & 64'hfe00707f; // @[Lookup.scala 31:38]
  wire  _T_19 = 64'h33 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_21 = 64'h1033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_23 = 64'h2033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_25 = 64'h3033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_27 = 64'h4033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_29 = 64'h5033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_31 = 64'h6033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_33 = 64'h7033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_35 = 64'h40000033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_37 = 64'h40005033 == _T_18; // @[Lookup.scala 31:38]
  wire [63:0] _T_38 = io_in_bits_instr & 64'h7f; // @[Lookup.scala 31:38]
  wire  _T_39 = 64'h17 == _T_38; // @[Lookup.scala 31:38]
  wire  _T_41 = 64'h37 == _T_38; // @[Lookup.scala 31:38]
  wire  _T_43 = 64'h6f == _T_38; // @[Lookup.scala 31:38]
  wire  _T_45 = 64'h67 == _T; // @[Lookup.scala 31:38]
  wire  _T_47 = 64'h63 == _T; // @[Lookup.scala 31:38]
  wire  _T_49 = 64'h1063 == _T; // @[Lookup.scala 31:38]
  wire  _T_51 = 64'h4063 == _T; // @[Lookup.scala 31:38]
  wire  _T_53 = 64'h5063 == _T; // @[Lookup.scala 31:38]
  wire  _T_55 = 64'h6063 == _T; // @[Lookup.scala 31:38]
  wire  _T_57 = 64'h7063 == _T; // @[Lookup.scala 31:38]
  wire  _T_59 = 64'h3 == _T; // @[Lookup.scala 31:38]
  wire  _T_61 = 64'h1003 == _T; // @[Lookup.scala 31:38]
  wire  _T_63 = 64'h2003 == _T; // @[Lookup.scala 31:38]
  wire  _T_65 = 64'h4003 == _T; // @[Lookup.scala 31:38]
  wire  _T_67 = 64'h5003 == _T; // @[Lookup.scala 31:38]
  wire  _T_69 = 64'h23 == _T; // @[Lookup.scala 31:38]
  wire  _T_71 = 64'h1023 == _T; // @[Lookup.scala 31:38]
  wire  _T_73 = 64'h2023 == _T; // @[Lookup.scala 31:38]
  wire  _T_75 = 64'h1b == _T; // @[Lookup.scala 31:38]
  wire  _T_77 = 64'h101b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_79 = 64'h501b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_81 = 64'h4000501b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_83 = 64'h103b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_85 = 64'h503b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_87 = 64'h4000503b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_89 = 64'h3b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_91 = 64'h4000003b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_93 = 64'h6003 == _T; // @[Lookup.scala 31:38]
  wire  _T_95 = 64'h3003 == _T; // @[Lookup.scala 31:38]
  wire  _T_97 = 64'h3023 == _T; // @[Lookup.scala 31:38]
  wire  _T_99 = 64'h6b == _T; // @[Lookup.scala 31:38]
  wire  _T_101 = 64'h2000033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_103 = 64'h2001033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_105 = 64'h2002033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_107 = 64'h2003033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_109 = 64'h2004033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_111 = 64'h2005033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_113 = 64'h2006033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_115 = 64'h2007033 == _T_18; // @[Lookup.scala 31:38]
  wire  _T_117 = 64'h200003b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_119 = 64'h200403b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_121 = 64'h200503b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_123 = 64'h200603b == _T_18; // @[Lookup.scala 31:38]
  wire  _T_125 = 64'h200703b == _T_18; // @[Lookup.scala 31:38]
  wire [63:0] _T_126 = io_in_bits_instr & 64'hffffffff; // @[Lookup.scala 31:38]
  wire  _T_127 = 64'h0 == _T_126; // @[Lookup.scala 31:38]
  wire [63:0] _T_128 = io_in_bits_instr & 64'he003; // @[Lookup.scala 31:38]
  wire  _T_129 = 64'h0 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_131 = 64'h4000 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_133 = 64'h6000 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_135 = 64'hc000 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_137 = 64'he000 == _T_128; // @[Lookup.scala 31:38]
  wire [63:0] _T_138 = io_in_bits_instr & 64'hef83; // @[Lookup.scala 31:38]
  wire  _T_139 = 64'h1 == _T_138; // @[Lookup.scala 31:38]
  wire  _T_141 = 64'h1 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_143 = 64'h2001 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_145 = 64'h4001 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_147 = 64'h6101 == _T_138; // @[Lookup.scala 31:38]
  wire  _T_149 = 64'h6001 == _T_128; // @[Lookup.scala 31:38]
  wire [63:0] _T_150 = io_in_bits_instr & 64'hec03; // @[Lookup.scala 31:38]
  wire  _T_151 = 64'h8001 == _T_150; // @[Lookup.scala 31:38]
  wire  _T_153 = 64'h8401 == _T_150; // @[Lookup.scala 31:38]
  wire  _T_155 = 64'h8801 == _T_150; // @[Lookup.scala 31:38]
  wire [63:0] _T_156 = io_in_bits_instr & 64'hfc63; // @[Lookup.scala 31:38]
  wire  _T_157 = 64'h8c01 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_159 = 64'h8c21 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_161 = 64'h8c41 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_163 = 64'h8c61 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_165 = 64'h9c01 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_167 = 64'h9c21 == _T_156; // @[Lookup.scala 31:38]
  wire  _T_169 = 64'ha001 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_171 = 64'hc001 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_173 = 64'he001 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_175 = 64'h2 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_177 = 64'h4002 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_179 = 64'h6002 == _T_128; // @[Lookup.scala 31:38]
  wire [63:0] _T_180 = io_in_bits_instr & 64'hf07f; // @[Lookup.scala 31:38]
  wire  _T_181 = 64'h8002 == _T_180; // @[Lookup.scala 31:38]
  wire [63:0] _T_182 = io_in_bits_instr & 64'hf003; // @[Lookup.scala 31:38]
  wire  _T_183 = 64'h8002 == _T_182; // @[Lookup.scala 31:38]
  wire [63:0] _T_184 = io_in_bits_instr & 64'hffff; // @[Lookup.scala 31:38]
  wire  _T_185 = 64'h9002 == _T_184; // @[Lookup.scala 31:38]
  wire  _T_187 = 64'h9002 == _T_180; // @[Lookup.scala 31:38]
  wire  _T_189 = 64'h9002 == _T_182; // @[Lookup.scala 31:38]
  wire  _T_191 = 64'hc002 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_193 = 64'he002 == _T_128; // @[Lookup.scala 31:38]
  wire  _T_195 = 64'h73 == _T_126; // @[Lookup.scala 31:38]
  wire  _T_197 = 64'h100073 == _T_126; // @[Lookup.scala 31:38]
  wire  _T_199 = 64'h30200073 == _T_126; // @[Lookup.scala 31:38]
  wire  _T_201 = 64'hf == _T; // @[Lookup.scala 31:38]
  wire  _T_203 = 64'h10500073 == _T_126; // @[Lookup.scala 31:38]
  wire  _T_205 = 64'h10200073 == _T_126; // @[Lookup.scala 31:38]
  wire [63:0] _T_206 = io_in_bits_instr & 64'hfe007fff; // @[Lookup.scala 31:38]
  wire  _T_207 = 64'h12000073 == _T_206; // @[Lookup.scala 31:38]
  wire [63:0] _T_208 = io_in_bits_instr & 64'hf9f0707f; // @[Lookup.scala 31:38]
  wire  _T_209 = 64'h1000302f == _T_208; // @[Lookup.scala 31:38]
  wire  _T_211 = 64'h1000202f == _T_208; // @[Lookup.scala 31:38]
  wire [63:0] _T_212 = io_in_bits_instr & 64'hf800707f; // @[Lookup.scala 31:38]
  wire  _T_213 = 64'h1800302f == _T_212; // @[Lookup.scala 31:38]
  wire  _T_215 = 64'h1800202f == _T_212; // @[Lookup.scala 31:38]
  wire [63:0] _T_216 = io_in_bits_instr & 64'hf800607f; // @[Lookup.scala 31:38]
  wire  _T_217 = 64'h800202f == _T_216; // @[Lookup.scala 31:38]
  wire  _T_219 = 64'h202f == _T_216; // @[Lookup.scala 31:38]
  wire  _T_221 = 64'h2000202f == _T_216; // @[Lookup.scala 31:38]
  wire  _T_223 = 64'h6000202f == _T_216; // @[Lookup.scala 31:38]
  wire  _T_225 = 64'h4000202f == _T_216; // @[Lookup.scala 31:38]
  wire  _T_227 = 64'h8000202f == _T_216; // @[Lookup.scala 31:38]
  wire  _T_229 = 64'ha000202f == _T_216; // @[Lookup.scala 31:38]
  wire  _T_231 = 64'hc000202f == _T_216; // @[Lookup.scala 31:38]
  wire  _T_233 = 64'he000202f == _T_216; // @[Lookup.scala 31:38]
  wire  _T_235 = 64'h1073 == _T; // @[Lookup.scala 31:38]
  wire  _T_237 = 64'h2073 == _T; // @[Lookup.scala 31:38]
  wire  _T_239 = 64'h3073 == _T; // @[Lookup.scala 31:38]
  wire  _T_241 = 64'h5073 == _T; // @[Lookup.scala 31:38]
  wire  _T_243 = 64'h6073 == _T; // @[Lookup.scala 31:38]
  wire  _T_245 = 64'h7073 == _T; // @[Lookup.scala 31:38]
  wire  _T_247 = 64'h100f == _T_126; // @[Lookup.scala 31:38]
  wire [2:0] _T_249 = _T_245 ? 3'h4 : {{2'd0}, _T_247}; // @[Lookup.scala 33:37]
  wire [2:0] _T_250 = _T_243 ? 3'h4 : _T_249; // @[Lookup.scala 33:37]
  wire [2:0] _T_251 = _T_241 ? 3'h4 : _T_250; // @[Lookup.scala 33:37]
  wire [2:0] _T_252 = _T_239 ? 3'h4 : _T_251; // @[Lookup.scala 33:37]
  wire [2:0] _T_253 = _T_237 ? 3'h4 : _T_252; // @[Lookup.scala 33:37]
  wire [2:0] _T_254 = _T_235 ? 3'h4 : _T_253; // @[Lookup.scala 33:37]
  wire [2:0] _T_255 = _T_233 ? 3'h5 : _T_254; // @[Lookup.scala 33:37]
  wire [2:0] _T_256 = _T_231 ? 3'h5 : _T_255; // @[Lookup.scala 33:37]
  wire [2:0] _T_257 = _T_229 ? 3'h5 : _T_256; // @[Lookup.scala 33:37]
  wire [2:0] _T_258 = _T_227 ? 3'h5 : _T_257; // @[Lookup.scala 33:37]
  wire [2:0] _T_259 = _T_225 ? 3'h5 : _T_258; // @[Lookup.scala 33:37]
  wire [2:0] _T_260 = _T_223 ? 3'h5 : _T_259; // @[Lookup.scala 33:37]
  wire [2:0] _T_261 = _T_221 ? 3'h5 : _T_260; // @[Lookup.scala 33:37]
  wire [2:0] _T_262 = _T_219 ? 3'h5 : _T_261; // @[Lookup.scala 33:37]
  wire [2:0] _T_263 = _T_217 ? 3'h5 : _T_262; // @[Lookup.scala 33:37]
  wire [3:0] _T_264 = _T_215 ? 4'hf : {{1'd0}, _T_263}; // @[Lookup.scala 33:37]
  wire [3:0] _T_265 = _T_213 ? 4'hf : _T_264; // @[Lookup.scala 33:37]
  wire [3:0] _T_266 = _T_211 ? 4'h4 : _T_265; // @[Lookup.scala 33:37]
  wire [3:0] _T_267 = _T_209 ? 4'h4 : _T_266; // @[Lookup.scala 33:37]
  wire [3:0] _T_268 = _T_207 ? 4'h5 : _T_267; // @[Lookup.scala 33:37]
  wire [3:0] _T_269 = _T_205 ? 4'h4 : _T_268; // @[Lookup.scala 33:37]
  wire [3:0] _T_270 = _T_203 ? 4'h4 : _T_269; // @[Lookup.scala 33:37]
  wire [3:0] _T_271 = _T_201 ? 4'h2 : _T_270; // @[Lookup.scala 33:37]
  wire [3:0] _T_272 = _T_199 ? 4'h4 : _T_271; // @[Lookup.scala 33:37]
  wire [3:0] _T_273 = _T_197 ? 4'h4 : _T_272; // @[Lookup.scala 33:37]
  wire [3:0] _T_274 = _T_195 ? 4'h4 : _T_273; // @[Lookup.scala 33:37]
  wire [3:0] _T_275 = _T_193 ? 4'h2 : _T_274; // @[Lookup.scala 33:37]
  wire [3:0] _T_276 = _T_191 ? 4'h2 : _T_275; // @[Lookup.scala 33:37]
  wire [3:0] _T_277 = _T_189 ? 4'h5 : _T_276; // @[Lookup.scala 33:37]
  wire [3:0] _T_278 = _T_187 ? 4'h4 : _T_277; // @[Lookup.scala 33:37]
  wire [3:0] _T_279 = _T_185 ? 4'h4 : _T_278; // @[Lookup.scala 33:37]
  wire [3:0] _T_280 = _T_183 ? 4'h5 : _T_279; // @[Lookup.scala 33:37]
  wire [3:0] _T_281 = _T_181 ? 4'h4 : _T_280; // @[Lookup.scala 33:37]
  wire [3:0] _T_282 = _T_179 ? 4'h4 : _T_281; // @[Lookup.scala 33:37]
  wire [3:0] _T_283 = _T_177 ? 4'h4 : _T_282; // @[Lookup.scala 33:37]
  wire [3:0] _T_284 = _T_175 ? 4'h4 : _T_283; // @[Lookup.scala 33:37]
  wire [3:0] _T_285 = _T_173 ? 4'h1 : _T_284; // @[Lookup.scala 33:37]
  wire [3:0] _T_286 = _T_171 ? 4'h1 : _T_285; // @[Lookup.scala 33:37]
  wire [3:0] _T_287 = _T_169 ? 4'h7 : _T_286; // @[Lookup.scala 33:37]
  wire [3:0] _T_288 = _T_167 ? 4'h5 : _T_287; // @[Lookup.scala 33:37]
  wire [3:0] _T_289 = _T_165 ? 4'h5 : _T_288; // @[Lookup.scala 33:37]
  wire [3:0] _T_290 = _T_163 ? 4'h5 : _T_289; // @[Lookup.scala 33:37]
  wire [3:0] _T_291 = _T_161 ? 4'h5 : _T_290; // @[Lookup.scala 33:37]
  wire [3:0] _T_292 = _T_159 ? 4'h5 : _T_291; // @[Lookup.scala 33:37]
  wire [3:0] _T_293 = _T_157 ? 4'h5 : _T_292; // @[Lookup.scala 33:37]
  wire [3:0] _T_294 = _T_155 ? 4'h4 : _T_293; // @[Lookup.scala 33:37]
  wire [3:0] _T_295 = _T_153 ? 4'h4 : _T_294; // @[Lookup.scala 33:37]
  wire [3:0] _T_296 = _T_151 ? 4'h4 : _T_295; // @[Lookup.scala 33:37]
  wire [3:0] _T_297 = _T_149 ? 4'h4 : _T_296; // @[Lookup.scala 33:37]
  wire [3:0] _T_298 = _T_147 ? 4'h4 : _T_297; // @[Lookup.scala 33:37]
  wire [3:0] _T_299 = _T_145 ? 4'h4 : _T_298; // @[Lookup.scala 33:37]
  wire [3:0] _T_300 = _T_143 ? 4'h4 : _T_299; // @[Lookup.scala 33:37]
  wire [3:0] _T_301 = _T_141 ? 4'h4 : _T_300; // @[Lookup.scala 33:37]
  wire [3:0] _T_302 = _T_139 ? 4'h4 : _T_301; // @[Lookup.scala 33:37]
  wire [3:0] _T_303 = _T_137 ? 4'h2 : _T_302; // @[Lookup.scala 33:37]
  wire [3:0] _T_304 = _T_135 ? 4'h2 : _T_303; // @[Lookup.scala 33:37]
  wire [3:0] _T_305 = _T_133 ? 4'h4 : _T_304; // @[Lookup.scala 33:37]
  wire [3:0] _T_306 = _T_131 ? 4'h4 : _T_305; // @[Lookup.scala 33:37]
  wire [3:0] _T_307 = _T_129 ? 4'h4 : _T_306; // @[Lookup.scala 33:37]
  wire [3:0] _T_308 = _T_127 ? 4'h0 : _T_307; // @[Lookup.scala 33:37]
  wire [3:0] _T_309 = _T_125 ? 4'h5 : _T_308; // @[Lookup.scala 33:37]
  wire [3:0] _T_310 = _T_123 ? 4'h5 : _T_309; // @[Lookup.scala 33:37]
  wire [3:0] _T_311 = _T_121 ? 4'h5 : _T_310; // @[Lookup.scala 33:37]
  wire [3:0] _T_312 = _T_119 ? 4'h5 : _T_311; // @[Lookup.scala 33:37]
  wire [3:0] _T_313 = _T_117 ? 4'h5 : _T_312; // @[Lookup.scala 33:37]
  wire [3:0] _T_314 = _T_115 ? 4'h5 : _T_313; // @[Lookup.scala 33:37]
  wire [3:0] _T_315 = _T_113 ? 4'h5 : _T_314; // @[Lookup.scala 33:37]
  wire [3:0] _T_316 = _T_111 ? 4'h5 : _T_315; // @[Lookup.scala 33:37]
  wire [3:0] _T_317 = _T_109 ? 4'h5 : _T_316; // @[Lookup.scala 33:37]
  wire [3:0] _T_318 = _T_107 ? 4'h5 : _T_317; // @[Lookup.scala 33:37]
  wire [3:0] _T_319 = _T_105 ? 4'h5 : _T_318; // @[Lookup.scala 33:37]
  wire [3:0] _T_320 = _T_103 ? 4'h5 : _T_319; // @[Lookup.scala 33:37]
  wire [3:0] _T_321 = _T_101 ? 4'h5 : _T_320; // @[Lookup.scala 33:37]
  wire [3:0] _T_322 = _T_99 ? 4'h4 : _T_321; // @[Lookup.scala 33:37]
  wire [3:0] _T_323 = _T_97 ? 4'h2 : _T_322; // @[Lookup.scala 33:37]
  wire [3:0] _T_324 = _T_95 ? 4'h4 : _T_323; // @[Lookup.scala 33:37]
  wire [3:0] _T_325 = _T_93 ? 4'h4 : _T_324; // @[Lookup.scala 33:37]
  wire [3:0] _T_326 = _T_91 ? 4'h5 : _T_325; // @[Lookup.scala 33:37]
  wire [3:0] _T_327 = _T_89 ? 4'h5 : _T_326; // @[Lookup.scala 33:37]
  wire [3:0] _T_328 = _T_87 ? 4'h5 : _T_327; // @[Lookup.scala 33:37]
  wire [3:0] _T_329 = _T_85 ? 4'h5 : _T_328; // @[Lookup.scala 33:37]
  wire [3:0] _T_330 = _T_83 ? 4'h5 : _T_329; // @[Lookup.scala 33:37]
  wire [3:0] _T_331 = _T_81 ? 4'h4 : _T_330; // @[Lookup.scala 33:37]
  wire [3:0] _T_332 = _T_79 ? 4'h4 : _T_331; // @[Lookup.scala 33:37]
  wire [3:0] _T_333 = _T_77 ? 4'h4 : _T_332; // @[Lookup.scala 33:37]
  wire [3:0] _T_334 = _T_75 ? 4'h4 : _T_333; // @[Lookup.scala 33:37]
  wire [3:0] _T_335 = _T_73 ? 4'h2 : _T_334; // @[Lookup.scala 33:37]
  wire [3:0] _T_336 = _T_71 ? 4'h2 : _T_335; // @[Lookup.scala 33:37]
  wire [3:0] _T_337 = _T_69 ? 4'h2 : _T_336; // @[Lookup.scala 33:37]
  wire [3:0] _T_338 = _T_67 ? 4'h4 : _T_337; // @[Lookup.scala 33:37]
  wire [3:0] _T_339 = _T_65 ? 4'h4 : _T_338; // @[Lookup.scala 33:37]
  wire [3:0] _T_340 = _T_63 ? 4'h4 : _T_339; // @[Lookup.scala 33:37]
  wire [3:0] _T_341 = _T_61 ? 4'h4 : _T_340; // @[Lookup.scala 33:37]
  wire [3:0] _T_342 = _T_59 ? 4'h4 : _T_341; // @[Lookup.scala 33:37]
  wire [3:0] _T_343 = _T_57 ? 4'h1 : _T_342; // @[Lookup.scala 33:37]
  wire [3:0] _T_344 = _T_55 ? 4'h1 : _T_343; // @[Lookup.scala 33:37]
  wire [3:0] _T_345 = _T_53 ? 4'h1 : _T_344; // @[Lookup.scala 33:37]
  wire [3:0] _T_346 = _T_51 ? 4'h1 : _T_345; // @[Lookup.scala 33:37]
  wire [3:0] _T_347 = _T_49 ? 4'h1 : _T_346; // @[Lookup.scala 33:37]
  wire [3:0] _T_348 = _T_47 ? 4'h1 : _T_347; // @[Lookup.scala 33:37]
  wire [3:0] _T_349 = _T_45 ? 4'h4 : _T_348; // @[Lookup.scala 33:37]
  wire [3:0] _T_350 = _T_43 ? 4'h7 : _T_349; // @[Lookup.scala 33:37]
  wire [3:0] _T_351 = _T_41 ? 4'h6 : _T_350; // @[Lookup.scala 33:37]
  wire [3:0] _T_352 = _T_39 ? 4'h6 : _T_351; // @[Lookup.scala 33:37]
  wire [3:0] _T_353 = _T_37 ? 4'h5 : _T_352; // @[Lookup.scala 33:37]
  wire [3:0] _T_354 = _T_35 ? 4'h5 : _T_353; // @[Lookup.scala 33:37]
  wire [3:0] _T_355 = _T_33 ? 4'h5 : _T_354; // @[Lookup.scala 33:37]
  wire [3:0] _T_356 = _T_31 ? 4'h5 : _T_355; // @[Lookup.scala 33:37]
  wire [3:0] _T_357 = _T_29 ? 4'h5 : _T_356; // @[Lookup.scala 33:37]
  wire [3:0] _T_358 = _T_27 ? 4'h5 : _T_357; // @[Lookup.scala 33:37]
  wire [3:0] _T_359 = _T_25 ? 4'h5 : _T_358; // @[Lookup.scala 33:37]
  wire [3:0] _T_360 = _T_23 ? 4'h5 : _T_359; // @[Lookup.scala 33:37]
  wire [3:0] _T_361 = _T_21 ? 4'h5 : _T_360; // @[Lookup.scala 33:37]
  wire [3:0] _T_362 = _T_19 ? 4'h5 : _T_361; // @[Lookup.scala 33:37]
  wire [3:0] _T_363 = _T_17 ? 4'h4 : _T_362; // @[Lookup.scala 33:37]
  wire [3:0] _T_364 = _T_15 ? 4'h4 : _T_363; // @[Lookup.scala 33:37]
  wire [3:0] _T_365 = _T_13 ? 4'h4 : _T_364; // @[Lookup.scala 33:37]
  wire [3:0] _T_366 = _T_11 ? 4'h4 : _T_365; // @[Lookup.scala 33:37]
  wire [3:0] _T_367 = _T_9 ? 4'h4 : _T_366; // @[Lookup.scala 33:37]
  wire [3:0] _T_368 = _T_7 ? 4'h4 : _T_367; // @[Lookup.scala 33:37]
  wire [3:0] _T_369 = _T_5 ? 4'h4 : _T_368; // @[Lookup.scala 33:37]
  wire [3:0] _T_370 = _T_3 ? 4'h4 : _T_369; // @[Lookup.scala 33:37]
  wire [3:0] decodeList_0 = _T_1 ? 4'h4 : _T_370; // @[Lookup.scala 33:37]
  wire [2:0] _T_371 = _T_247 ? 3'h4 : 3'h3; // @[Lookup.scala 33:37]
  wire [2:0] _T_372 = _T_245 ? 3'h3 : _T_371; // @[Lookup.scala 33:37]
  wire [2:0] _T_373 = _T_243 ? 3'h3 : _T_372; // @[Lookup.scala 33:37]
  wire [2:0] _T_374 = _T_241 ? 3'h3 : _T_373; // @[Lookup.scala 33:37]
  wire [2:0] _T_375 = _T_239 ? 3'h3 : _T_374; // @[Lookup.scala 33:37]
  wire [2:0] _T_376 = _T_237 ? 3'h3 : _T_375; // @[Lookup.scala 33:37]
  wire [2:0] _T_377 = _T_235 ? 3'h3 : _T_376; // @[Lookup.scala 33:37]
  wire [2:0] _T_378 = _T_233 ? 3'h1 : _T_377; // @[Lookup.scala 33:37]
  wire [2:0] _T_379 = _T_231 ? 3'h1 : _T_378; // @[Lookup.scala 33:37]
  wire [2:0] _T_380 = _T_229 ? 3'h1 : _T_379; // @[Lookup.scala 33:37]
  wire [2:0] _T_381 = _T_227 ? 3'h1 : _T_380; // @[Lookup.scala 33:37]
  wire [2:0] _T_382 = _T_225 ? 3'h1 : _T_381; // @[Lookup.scala 33:37]
  wire [2:0] _T_383 = _T_223 ? 3'h1 : _T_382; // @[Lookup.scala 33:37]
  wire [2:0] _T_384 = _T_221 ? 3'h1 : _T_383; // @[Lookup.scala 33:37]
  wire [2:0] _T_385 = _T_219 ? 3'h1 : _T_384; // @[Lookup.scala 33:37]
  wire [2:0] _T_386 = _T_217 ? 3'h1 : _T_385; // @[Lookup.scala 33:37]
  wire [2:0] _T_387 = _T_215 ? 3'h1 : _T_386; // @[Lookup.scala 33:37]
  wire [2:0] _T_388 = _T_213 ? 3'h1 : _T_387; // @[Lookup.scala 33:37]
  wire [2:0] _T_389 = _T_211 ? 3'h1 : _T_388; // @[Lookup.scala 33:37]
  wire [2:0] _T_390 = _T_209 ? 3'h1 : _T_389; // @[Lookup.scala 33:37]
  wire [2:0] _T_391 = _T_207 ? 3'h4 : _T_390; // @[Lookup.scala 33:37]
  wire [2:0] _T_392 = _T_205 ? 3'h3 : _T_391; // @[Lookup.scala 33:37]
  wire [2:0] _T_393 = _T_203 ? 3'h0 : _T_392; // @[Lookup.scala 33:37]
  wire [2:0] _T_394 = _T_201 ? 3'h4 : _T_393; // @[Lookup.scala 33:37]
  wire [2:0] _T_395 = _T_199 ? 3'h3 : _T_394; // @[Lookup.scala 33:37]
  wire [2:0] _T_396 = _T_197 ? 3'h3 : _T_395; // @[Lookup.scala 33:37]
  wire [2:0] _T_397 = _T_195 ? 3'h3 : _T_396; // @[Lookup.scala 33:37]
  wire [2:0] _T_398 = _T_193 ? 3'h1 : _T_397; // @[Lookup.scala 33:37]
  wire [2:0] _T_399 = _T_191 ? 3'h1 : _T_398; // @[Lookup.scala 33:37]
  wire [2:0] _T_400 = _T_189 ? 3'h0 : _T_399; // @[Lookup.scala 33:37]
  wire [2:0] _T_401 = _T_187 ? 3'h0 : _T_400; // @[Lookup.scala 33:37]
  wire [2:0] _T_402 = _T_185 ? 3'h3 : _T_401; // @[Lookup.scala 33:37]
  wire [2:0] _T_403 = _T_183 ? 3'h0 : _T_402; // @[Lookup.scala 33:37]
  wire [2:0] _T_404 = _T_181 ? 3'h0 : _T_403; // @[Lookup.scala 33:37]
  wire [2:0] _T_405 = _T_179 ? 3'h1 : _T_404; // @[Lookup.scala 33:37]
  wire [2:0] _T_406 = _T_177 ? 3'h1 : _T_405; // @[Lookup.scala 33:37]
  wire [2:0] _T_407 = _T_175 ? 3'h0 : _T_406; // @[Lookup.scala 33:37]
  wire [2:0] _T_408 = _T_173 ? 3'h0 : _T_407; // @[Lookup.scala 33:37]
  wire [2:0] _T_409 = _T_171 ? 3'h0 : _T_408; // @[Lookup.scala 33:37]
  wire [2:0] _T_410 = _T_169 ? 3'h0 : _T_409; // @[Lookup.scala 33:37]
  wire [2:0] _T_411 = _T_167 ? 3'h0 : _T_410; // @[Lookup.scala 33:37]
  wire [2:0] _T_412 = _T_165 ? 3'h0 : _T_411; // @[Lookup.scala 33:37]
  wire [2:0] _T_413 = _T_163 ? 3'h0 : _T_412; // @[Lookup.scala 33:37]
  wire [2:0] _T_414 = _T_161 ? 3'h0 : _T_413; // @[Lookup.scala 33:37]
  wire [2:0] _T_415 = _T_159 ? 3'h0 : _T_414; // @[Lookup.scala 33:37]
  wire [2:0] _T_416 = _T_157 ? 3'h0 : _T_415; // @[Lookup.scala 33:37]
  wire [2:0] _T_417 = _T_155 ? 3'h0 : _T_416; // @[Lookup.scala 33:37]
  wire [2:0] _T_418 = _T_153 ? 3'h0 : _T_417; // @[Lookup.scala 33:37]
  wire [2:0] _T_419 = _T_151 ? 3'h0 : _T_418; // @[Lookup.scala 33:37]
  wire [2:0] _T_420 = _T_149 ? 3'h0 : _T_419; // @[Lookup.scala 33:37]
  wire [2:0] _T_421 = _T_147 ? 3'h0 : _T_420; // @[Lookup.scala 33:37]
  wire [2:0] _T_422 = _T_145 ? 3'h0 : _T_421; // @[Lookup.scala 33:37]
  wire [2:0] _T_423 = _T_143 ? 3'h0 : _T_422; // @[Lookup.scala 33:37]
  wire [2:0] _T_424 = _T_141 ? 3'h0 : _T_423; // @[Lookup.scala 33:37]
  wire [2:0] _T_425 = _T_139 ? 3'h0 : _T_424; // @[Lookup.scala 33:37]
  wire [2:0] _T_426 = _T_137 ? 3'h1 : _T_425; // @[Lookup.scala 33:37]
  wire [2:0] _T_427 = _T_135 ? 3'h1 : _T_426; // @[Lookup.scala 33:37]
  wire [2:0] _T_428 = _T_133 ? 3'h1 : _T_427; // @[Lookup.scala 33:37]
  wire [2:0] _T_429 = _T_131 ? 3'h1 : _T_428; // @[Lookup.scala 33:37]
  wire [2:0] _T_430 = _T_129 ? 3'h0 : _T_429; // @[Lookup.scala 33:37]
  wire [2:0] _T_431 = _T_127 ? 3'h3 : _T_430; // @[Lookup.scala 33:37]
  wire [2:0] _T_432 = _T_125 ? 3'h2 : _T_431; // @[Lookup.scala 33:37]
  wire [2:0] _T_433 = _T_123 ? 3'h2 : _T_432; // @[Lookup.scala 33:37]
  wire [2:0] _T_434 = _T_121 ? 3'h2 : _T_433; // @[Lookup.scala 33:37]
  wire [2:0] _T_435 = _T_119 ? 3'h2 : _T_434; // @[Lookup.scala 33:37]
  wire [2:0] _T_436 = _T_117 ? 3'h2 : _T_435; // @[Lookup.scala 33:37]
  wire [2:0] _T_437 = _T_115 ? 3'h2 : _T_436; // @[Lookup.scala 33:37]
  wire [2:0] _T_438 = _T_113 ? 3'h2 : _T_437; // @[Lookup.scala 33:37]
  wire [2:0] _T_439 = _T_111 ? 3'h2 : _T_438; // @[Lookup.scala 33:37]
  wire [2:0] _T_440 = _T_109 ? 3'h2 : _T_439; // @[Lookup.scala 33:37]
  wire [2:0] _T_441 = _T_107 ? 3'h2 : _T_440; // @[Lookup.scala 33:37]
  wire [2:0] _T_442 = _T_105 ? 3'h2 : _T_441; // @[Lookup.scala 33:37]
  wire [2:0] _T_443 = _T_103 ? 3'h2 : _T_442; // @[Lookup.scala 33:37]
  wire [2:0] _T_444 = _T_101 ? 3'h2 : _T_443; // @[Lookup.scala 33:37]
  wire [2:0] _T_445 = _T_99 ? 3'h3 : _T_444; // @[Lookup.scala 33:37]
  wire [2:0] _T_446 = _T_97 ? 3'h1 : _T_445; // @[Lookup.scala 33:37]
  wire [2:0] _T_447 = _T_95 ? 3'h1 : _T_446; // @[Lookup.scala 33:37]
  wire [2:0] _T_448 = _T_93 ? 3'h1 : _T_447; // @[Lookup.scala 33:37]
  wire [2:0] _T_449 = _T_91 ? 3'h0 : _T_448; // @[Lookup.scala 33:37]
  wire [2:0] _T_450 = _T_89 ? 3'h0 : _T_449; // @[Lookup.scala 33:37]
  wire [2:0] _T_451 = _T_87 ? 3'h0 : _T_450; // @[Lookup.scala 33:37]
  wire [2:0] _T_452 = _T_85 ? 3'h0 : _T_451; // @[Lookup.scala 33:37]
  wire [2:0] _T_453 = _T_83 ? 3'h0 : _T_452; // @[Lookup.scala 33:37]
  wire [2:0] _T_454 = _T_81 ? 3'h0 : _T_453; // @[Lookup.scala 33:37]
  wire [2:0] _T_455 = _T_79 ? 3'h0 : _T_454; // @[Lookup.scala 33:37]
  wire [2:0] _T_456 = _T_77 ? 3'h0 : _T_455; // @[Lookup.scala 33:37]
  wire [2:0] _T_457 = _T_75 ? 3'h0 : _T_456; // @[Lookup.scala 33:37]
  wire [2:0] _T_458 = _T_73 ? 3'h1 : _T_457; // @[Lookup.scala 33:37]
  wire [2:0] _T_459 = _T_71 ? 3'h1 : _T_458; // @[Lookup.scala 33:37]
  wire [2:0] _T_460 = _T_69 ? 3'h1 : _T_459; // @[Lookup.scala 33:37]
  wire [2:0] _T_461 = _T_67 ? 3'h1 : _T_460; // @[Lookup.scala 33:37]
  wire [2:0] _T_462 = _T_65 ? 3'h1 : _T_461; // @[Lookup.scala 33:37]
  wire [2:0] _T_463 = _T_63 ? 3'h1 : _T_462; // @[Lookup.scala 33:37]
  wire [2:0] _T_464 = _T_61 ? 3'h1 : _T_463; // @[Lookup.scala 33:37]
  wire [2:0] _T_465 = _T_59 ? 3'h1 : _T_464; // @[Lookup.scala 33:37]
  wire [2:0] _T_466 = _T_57 ? 3'h0 : _T_465; // @[Lookup.scala 33:37]
  wire [2:0] _T_467 = _T_55 ? 3'h0 : _T_466; // @[Lookup.scala 33:37]
  wire [2:0] _T_468 = _T_53 ? 3'h0 : _T_467; // @[Lookup.scala 33:37]
  wire [2:0] _T_469 = _T_51 ? 3'h0 : _T_468; // @[Lookup.scala 33:37]
  wire [2:0] _T_470 = _T_49 ? 3'h0 : _T_469; // @[Lookup.scala 33:37]
  wire [2:0] _T_471 = _T_47 ? 3'h0 : _T_470; // @[Lookup.scala 33:37]
  wire [2:0] _T_472 = _T_45 ? 3'h0 : _T_471; // @[Lookup.scala 33:37]
  wire [2:0] _T_473 = _T_43 ? 3'h0 : _T_472; // @[Lookup.scala 33:37]
  wire [2:0] _T_474 = _T_41 ? 3'h0 : _T_473; // @[Lookup.scala 33:37]
  wire [2:0] _T_475 = _T_39 ? 3'h0 : _T_474; // @[Lookup.scala 33:37]
  wire [2:0] _T_476 = _T_37 ? 3'h0 : _T_475; // @[Lookup.scala 33:37]
  wire [2:0] _T_477 = _T_35 ? 3'h0 : _T_476; // @[Lookup.scala 33:37]
  wire [2:0] _T_478 = _T_33 ? 3'h0 : _T_477; // @[Lookup.scala 33:37]
  wire [2:0] _T_479 = _T_31 ? 3'h0 : _T_478; // @[Lookup.scala 33:37]
  wire [2:0] _T_480 = _T_29 ? 3'h0 : _T_479; // @[Lookup.scala 33:37]
  wire [2:0] _T_481 = _T_27 ? 3'h0 : _T_480; // @[Lookup.scala 33:37]
  wire [2:0] _T_482 = _T_25 ? 3'h0 : _T_481; // @[Lookup.scala 33:37]
  wire [2:0] _T_483 = _T_23 ? 3'h0 : _T_482; // @[Lookup.scala 33:37]
  wire [2:0] _T_484 = _T_21 ? 3'h0 : _T_483; // @[Lookup.scala 33:37]
  wire [2:0] _T_485 = _T_19 ? 3'h0 : _T_484; // @[Lookup.scala 33:37]
  wire [2:0] _T_486 = _T_17 ? 3'h0 : _T_485; // @[Lookup.scala 33:37]
  wire [2:0] _T_487 = _T_15 ? 3'h0 : _T_486; // @[Lookup.scala 33:37]
  wire [2:0] _T_488 = _T_13 ? 3'h0 : _T_487; // @[Lookup.scala 33:37]
  wire [2:0] _T_489 = _T_11 ? 3'h0 : _T_488; // @[Lookup.scala 33:37]
  wire [2:0] _T_490 = _T_9 ? 3'h0 : _T_489; // @[Lookup.scala 33:37]
  wire [2:0] _T_491 = _T_7 ? 3'h0 : _T_490; // @[Lookup.scala 33:37]
  wire [2:0] _T_492 = _T_5 ? 3'h0 : _T_491; // @[Lookup.scala 33:37]
  wire [2:0] _T_493 = _T_3 ? 3'h0 : _T_492; // @[Lookup.scala 33:37]
  wire [2:0] decodeList_1 = _T_1 ? 3'h0 : _T_493; // @[Lookup.scala 33:37]
  wire [2:0] _T_495 = _T_245 ? 3'h7 : {{2'd0}, _T_247}; // @[Lookup.scala 33:37]
  wire [2:0] _T_496 = _T_243 ? 3'h6 : _T_495; // @[Lookup.scala 33:37]
  wire [2:0] _T_497 = _T_241 ? 3'h5 : _T_496; // @[Lookup.scala 33:37]
  wire [2:0] _T_498 = _T_239 ? 3'h3 : _T_497; // @[Lookup.scala 33:37]
  wire [2:0] _T_499 = _T_237 ? 3'h2 : _T_498; // @[Lookup.scala 33:37]
  wire [2:0] _T_500 = _T_235 ? 3'h1 : _T_499; // @[Lookup.scala 33:37]
  wire [5:0] _T_501 = _T_233 ? 6'h32 : {{3'd0}, _T_500}; // @[Lookup.scala 33:37]
  wire [5:0] _T_502 = _T_231 ? 6'h31 : _T_501; // @[Lookup.scala 33:37]
  wire [5:0] _T_503 = _T_229 ? 6'h30 : _T_502; // @[Lookup.scala 33:37]
  wire [5:0] _T_504 = _T_227 ? 6'h37 : _T_503; // @[Lookup.scala 33:37]
  wire [5:0] _T_505 = _T_225 ? 6'h26 : _T_504; // @[Lookup.scala 33:37]
  wire [5:0] _T_506 = _T_223 ? 6'h25 : _T_505; // @[Lookup.scala 33:37]
  wire [5:0] _T_507 = _T_221 ? 6'h24 : _T_506; // @[Lookup.scala 33:37]
  wire [6:0] _T_508 = _T_219 ? 7'h63 : {{1'd0}, _T_507}; // @[Lookup.scala 33:37]
  wire [6:0] _T_509 = _T_217 ? 7'h22 : _T_508; // @[Lookup.scala 33:37]
  wire [6:0] _T_510 = _T_215 ? 7'h21 : _T_509; // @[Lookup.scala 33:37]
  wire [6:0] _T_511 = _T_213 ? 7'h21 : _T_510; // @[Lookup.scala 33:37]
  wire [6:0] _T_512 = _T_211 ? 7'h20 : _T_511; // @[Lookup.scala 33:37]
  wire [6:0] _T_513 = _T_209 ? 7'h20 : _T_512; // @[Lookup.scala 33:37]
  wire [6:0] _T_514 = _T_207 ? 7'h2 : _T_513; // @[Lookup.scala 33:37]
  wire [6:0] _T_515 = _T_205 ? 7'h0 : _T_514; // @[Lookup.scala 33:37]
  wire [6:0] _T_516 = _T_203 ? 7'h40 : _T_515; // @[Lookup.scala 33:37]
  wire [6:0] _T_517 = _T_201 ? 7'h0 : _T_516; // @[Lookup.scala 33:37]
  wire [6:0] _T_518 = _T_199 ? 7'h0 : _T_517; // @[Lookup.scala 33:37]
  wire [6:0] _T_519 = _T_197 ? 7'h0 : _T_518; // @[Lookup.scala 33:37]
  wire [6:0] _T_520 = _T_195 ? 7'h0 : _T_519; // @[Lookup.scala 33:37]
  wire [6:0] _T_521 = _T_193 ? 7'hb : _T_520; // @[Lookup.scala 33:37]
  wire [6:0] _T_522 = _T_191 ? 7'ha : _T_521; // @[Lookup.scala 33:37]
  wire [6:0] _T_523 = _T_189 ? 7'h40 : _T_522; // @[Lookup.scala 33:37]
  wire [6:0] _T_524 = _T_187 ? 7'h5a : _T_523; // @[Lookup.scala 33:37]
  wire [6:0] _T_525 = _T_185 ? 7'h0 : _T_524; // @[Lookup.scala 33:37]
  wire [6:0] _T_526 = _T_183 ? 7'h40 : _T_525; // @[Lookup.scala 33:37]
  wire [6:0] _T_527 = _T_181 ? 7'h5a : _T_526; // @[Lookup.scala 33:37]
  wire [6:0] _T_528 = _T_179 ? 7'h3 : _T_527; // @[Lookup.scala 33:37]
  wire [6:0] _T_529 = _T_177 ? 7'h2 : _T_528; // @[Lookup.scala 33:37]
  wire [6:0] _T_530 = _T_175 ? 7'h1 : _T_529; // @[Lookup.scala 33:37]
  wire [6:0] _T_531 = _T_173 ? 7'h11 : _T_530; // @[Lookup.scala 33:37]
  wire [6:0] _T_532 = _T_171 ? 7'h10 : _T_531; // @[Lookup.scala 33:37]
  wire [6:0] _T_533 = _T_169 ? 7'h58 : _T_532; // @[Lookup.scala 33:37]
  wire [6:0] _T_534 = _T_167 ? 7'h60 : _T_533; // @[Lookup.scala 33:37]
  wire [6:0] _T_535 = _T_165 ? 7'h28 : _T_534; // @[Lookup.scala 33:37]
  wire [6:0] _T_536 = _T_163 ? 7'h7 : _T_535; // @[Lookup.scala 33:37]
  wire [6:0] _T_537 = _T_161 ? 7'h6 : _T_536; // @[Lookup.scala 33:37]
  wire [6:0] _T_538 = _T_159 ? 7'h4 : _T_537; // @[Lookup.scala 33:37]
  wire [6:0] _T_539 = _T_157 ? 7'h8 : _T_538; // @[Lookup.scala 33:37]
  wire [6:0] _T_540 = _T_155 ? 7'h7 : _T_539; // @[Lookup.scala 33:37]
  wire [6:0] _T_541 = _T_153 ? 7'hd : _T_540; // @[Lookup.scala 33:37]
  wire [6:0] _T_542 = _T_151 ? 7'h5 : _T_541; // @[Lookup.scala 33:37]
  wire [6:0] _T_543 = _T_149 ? 7'h40 : _T_542; // @[Lookup.scala 33:37]
  wire [6:0] _T_544 = _T_147 ? 7'h40 : _T_543; // @[Lookup.scala 33:37]
  wire [6:0] _T_545 = _T_145 ? 7'h40 : _T_544; // @[Lookup.scala 33:37]
  wire [6:0] _T_546 = _T_143 ? 7'h60 : _T_545; // @[Lookup.scala 33:37]
  wire [6:0] _T_547 = _T_141 ? 7'h40 : _T_546; // @[Lookup.scala 33:37]
  wire [6:0] _T_548 = _T_139 ? 7'h40 : _T_547; // @[Lookup.scala 33:37]
  wire [6:0] _T_549 = _T_137 ? 7'hb : _T_548; // @[Lookup.scala 33:37]
  wire [6:0] _T_550 = _T_135 ? 7'ha : _T_549; // @[Lookup.scala 33:37]
  wire [6:0] _T_551 = _T_133 ? 7'h3 : _T_550; // @[Lookup.scala 33:37]
  wire [6:0] _T_552 = _T_131 ? 7'h2 : _T_551; // @[Lookup.scala 33:37]
  wire [6:0] _T_553 = _T_129 ? 7'h40 : _T_552; // @[Lookup.scala 33:37]
  wire [6:0] _T_554 = _T_127 ? 7'h0 : _T_553; // @[Lookup.scala 33:37]
  wire [6:0] _T_555 = _T_125 ? 7'hf : _T_554; // @[Lookup.scala 33:37]
  wire [6:0] _T_556 = _T_123 ? 7'he : _T_555; // @[Lookup.scala 33:37]
  wire [6:0] _T_557 = _T_121 ? 7'hd : _T_556; // @[Lookup.scala 33:37]
  wire [6:0] _T_558 = _T_119 ? 7'hc : _T_557; // @[Lookup.scala 33:37]
  wire [6:0] _T_559 = _T_117 ? 7'h8 : _T_558; // @[Lookup.scala 33:37]
  wire [6:0] _T_560 = _T_115 ? 7'h7 : _T_559; // @[Lookup.scala 33:37]
  wire [6:0] _T_561 = _T_113 ? 7'h6 : _T_560; // @[Lookup.scala 33:37]
  wire [6:0] _T_562 = _T_111 ? 7'h5 : _T_561; // @[Lookup.scala 33:37]
  wire [6:0] _T_563 = _T_109 ? 7'h4 : _T_562; // @[Lookup.scala 33:37]
  wire [6:0] _T_564 = _T_107 ? 7'h3 : _T_563; // @[Lookup.scala 33:37]
  wire [6:0] _T_565 = _T_105 ? 7'h2 : _T_564; // @[Lookup.scala 33:37]
  wire [6:0] _T_566 = _T_103 ? 7'h1 : _T_565; // @[Lookup.scala 33:37]
  wire [6:0] _T_567 = _T_101 ? 7'h0 : _T_566; // @[Lookup.scala 33:37]
  wire [6:0] _T_568 = _T_99 ? 7'h2 : _T_567; // @[Lookup.scala 33:37]
  wire [6:0] _T_569 = _T_97 ? 7'hb : _T_568; // @[Lookup.scala 33:37]
  wire [6:0] _T_570 = _T_95 ? 7'h3 : _T_569; // @[Lookup.scala 33:37]
  wire [6:0] _T_571 = _T_93 ? 7'h6 : _T_570; // @[Lookup.scala 33:37]
  wire [6:0] _T_572 = _T_91 ? 7'h28 : _T_571; // @[Lookup.scala 33:37]
  wire [6:0] _T_573 = _T_89 ? 7'h60 : _T_572; // @[Lookup.scala 33:37]
  wire [6:0] _T_574 = _T_87 ? 7'h2d : _T_573; // @[Lookup.scala 33:37]
  wire [6:0] _T_575 = _T_85 ? 7'h25 : _T_574; // @[Lookup.scala 33:37]
  wire [6:0] _T_576 = _T_83 ? 7'h21 : _T_575; // @[Lookup.scala 33:37]
  wire [6:0] _T_577 = _T_81 ? 7'h2d : _T_576; // @[Lookup.scala 33:37]
  wire [6:0] _T_578 = _T_79 ? 7'h25 : _T_577; // @[Lookup.scala 33:37]
  wire [6:0] _T_579 = _T_77 ? 7'h21 : _T_578; // @[Lookup.scala 33:37]
  wire [6:0] _T_580 = _T_75 ? 7'h60 : _T_579; // @[Lookup.scala 33:37]
  wire [6:0] _T_581 = _T_73 ? 7'ha : _T_580; // @[Lookup.scala 33:37]
  wire [6:0] _T_582 = _T_71 ? 7'h9 : _T_581; // @[Lookup.scala 33:37]
  wire [6:0] _T_583 = _T_69 ? 7'h8 : _T_582; // @[Lookup.scala 33:37]
  wire [6:0] _T_584 = _T_67 ? 7'h5 : _T_583; // @[Lookup.scala 33:37]
  wire [6:0] _T_585 = _T_65 ? 7'h4 : _T_584; // @[Lookup.scala 33:37]
  wire [6:0] _T_586 = _T_63 ? 7'h2 : _T_585; // @[Lookup.scala 33:37]
  wire [6:0] _T_587 = _T_61 ? 7'h1 : _T_586; // @[Lookup.scala 33:37]
  wire [6:0] _T_588 = _T_59 ? 7'h0 : _T_587; // @[Lookup.scala 33:37]
  wire [6:0] _T_589 = _T_57 ? 7'h17 : _T_588; // @[Lookup.scala 33:37]
  wire [6:0] _T_590 = _T_55 ? 7'h16 : _T_589; // @[Lookup.scala 33:37]
  wire [6:0] _T_591 = _T_53 ? 7'h15 : _T_590; // @[Lookup.scala 33:37]
  wire [6:0] _T_592 = _T_51 ? 7'h14 : _T_591; // @[Lookup.scala 33:37]
  wire [6:0] _T_593 = _T_49 ? 7'h11 : _T_592; // @[Lookup.scala 33:37]
  wire [6:0] _T_594 = _T_47 ? 7'h10 : _T_593; // @[Lookup.scala 33:37]
  wire [6:0] _T_595 = _T_45 ? 7'h5a : _T_594; // @[Lookup.scala 33:37]
  wire [6:0] _T_596 = _T_43 ? 7'h58 : _T_595; // @[Lookup.scala 33:37]
  wire [6:0] _T_597 = _T_41 ? 7'h40 : _T_596; // @[Lookup.scala 33:37]
  wire [6:0] _T_598 = _T_39 ? 7'h40 : _T_597; // @[Lookup.scala 33:37]
  wire [6:0] _T_599 = _T_37 ? 7'hd : _T_598; // @[Lookup.scala 33:37]
  wire [6:0] _T_600 = _T_35 ? 7'h8 : _T_599; // @[Lookup.scala 33:37]
  wire [6:0] _T_601 = _T_33 ? 7'h7 : _T_600; // @[Lookup.scala 33:37]
  wire [6:0] _T_602 = _T_31 ? 7'h6 : _T_601; // @[Lookup.scala 33:37]
  wire [6:0] _T_603 = _T_29 ? 7'h5 : _T_602; // @[Lookup.scala 33:37]
  wire [6:0] _T_604 = _T_27 ? 7'h4 : _T_603; // @[Lookup.scala 33:37]
  wire [6:0] _T_605 = _T_25 ? 7'h3 : _T_604; // @[Lookup.scala 33:37]
  wire [6:0] _T_606 = _T_23 ? 7'h2 : _T_605; // @[Lookup.scala 33:37]
  wire [6:0] _T_607 = _T_21 ? 7'h1 : _T_606; // @[Lookup.scala 33:37]
  wire [6:0] _T_608 = _T_19 ? 7'h40 : _T_607; // @[Lookup.scala 33:37]
  wire [6:0] _T_609 = _T_17 ? 7'hd : _T_608; // @[Lookup.scala 33:37]
  wire [6:0] _T_610 = _T_15 ? 7'h7 : _T_609; // @[Lookup.scala 33:37]
  wire [6:0] _T_611 = _T_13 ? 7'h6 : _T_610; // @[Lookup.scala 33:37]
  wire [6:0] _T_612 = _T_11 ? 7'h5 : _T_611; // @[Lookup.scala 33:37]
  wire [6:0] _T_613 = _T_9 ? 7'h4 : _T_612; // @[Lookup.scala 33:37]
  wire [6:0] _T_614 = _T_7 ? 7'h3 : _T_613; // @[Lookup.scala 33:37]
  wire [6:0] _T_615 = _T_5 ? 7'h2 : _T_614; // @[Lookup.scala 33:37]
  wire [6:0] _T_616 = _T_3 ? 7'h1 : _T_615; // @[Lookup.scala 33:37]
  wire [6:0] decodeList_2 = _T_1 ? 7'h40 : _T_616; // @[Lookup.scala 33:37]
  wire  hasIntr = |intrVecIDU; // @[IDU.scala 170:22]
  wire  _T_617 = hasIntr | io_in_bits_exceptionVec_12; // @[IDU.scala 36:84]
  wire  _T_618 = _T_617 | io_out_bits_cf_exceptionVec_1; // @[IDU.scala 36:127]
  wire [3:0] instrType = _T_618 ? 4'h0 : decodeList_0; // @[IDU.scala 36:75]
  wire [2:0] fuType = _T_618 ? 3'h3 : decodeList_1; // @[IDU.scala 36:75]
  wire [6:0] fuOpType = _T_618 ? 7'h0 : decodeList_2; // @[IDU.scala 36:75]
  wire  isRVC = io_in_bits_instr[1:0] != 2'h3; // @[IDU.scala 38:45]
  wire [4:0] _T_690 = _T_193 ? 5'h3 : 5'h10; // @[Lookup.scala 33:37]
  wire [4:0] _T_691 = _T_191 ? 5'h2 : _T_690; // @[Lookup.scala 33:37]
  wire [4:0] _T_692 = _T_189 ? 5'h10 : _T_691; // @[Lookup.scala 33:37]
  wire [4:0] _T_693 = _T_187 ? 5'h10 : _T_692; // @[Lookup.scala 33:37]
  wire [4:0] _T_694 = _T_185 ? 5'hf : _T_693; // @[Lookup.scala 33:37]
  wire [4:0] _T_695 = _T_183 ? 5'h10 : _T_694; // @[Lookup.scala 33:37]
  wire [4:0] _T_696 = _T_181 ? 5'h10 : _T_695; // @[Lookup.scala 33:37]
  wire [4:0] _T_697 = _T_179 ? 5'h1 : _T_696; // @[Lookup.scala 33:37]
  wire [4:0] _T_698 = _T_177 ? 5'h0 : _T_697; // @[Lookup.scala 33:37]
  wire [4:0] _T_699 = _T_175 ? 5'ha : _T_698; // @[Lookup.scala 33:37]
  wire [4:0] _T_700 = _T_173 ? 5'h9 : _T_699; // @[Lookup.scala 33:37]
  wire [4:0] _T_701 = _T_171 ? 5'h9 : _T_700; // @[Lookup.scala 33:37]
  wire [4:0] _T_702 = _T_169 ? 5'h8 : _T_701; // @[Lookup.scala 33:37]
  wire [4:0] _T_703 = _T_167 ? 5'h10 : _T_702; // @[Lookup.scala 33:37]
  wire [4:0] _T_704 = _T_165 ? 5'h10 : _T_703; // @[Lookup.scala 33:37]
  wire [4:0] _T_705 = _T_163 ? 5'h10 : _T_704; // @[Lookup.scala 33:37]
  wire [4:0] _T_706 = _T_161 ? 5'h10 : _T_705; // @[Lookup.scala 33:37]
  wire [4:0] _T_707 = _T_159 ? 5'h10 : _T_706; // @[Lookup.scala 33:37]
  wire [4:0] _T_708 = _T_157 ? 5'h10 : _T_707; // @[Lookup.scala 33:37]
  wire [4:0] _T_709 = _T_155 ? 5'ha : _T_708; // @[Lookup.scala 33:37]
  wire [4:0] _T_710 = _T_153 ? 5'ha : _T_709; // @[Lookup.scala 33:37]
  wire [4:0] _T_711 = _T_151 ? 5'ha : _T_710; // @[Lookup.scala 33:37]
  wire [4:0] _T_712 = _T_149 ? 5'hb : _T_711; // @[Lookup.scala 33:37]
  wire [4:0] _T_713 = _T_147 ? 5'hd : _T_712; // @[Lookup.scala 33:37]
  wire [4:0] _T_714 = _T_145 ? 5'ha : _T_713; // @[Lookup.scala 33:37]
  wire [4:0] _T_715 = _T_143 ? 5'hc : _T_714; // @[Lookup.scala 33:37]
  wire [4:0] _T_716 = _T_141 ? 5'hc : _T_715; // @[Lookup.scala 33:37]
  wire [4:0] _T_717 = _T_139 ? 5'h10 : _T_716; // @[Lookup.scala 33:37]
  wire [4:0] _T_718 = _T_137 ? 5'h5 : _T_717; // @[Lookup.scala 33:37]
  wire [4:0] _T_719 = _T_135 ? 5'h4 : _T_718; // @[Lookup.scala 33:37]
  wire [4:0] _T_720 = _T_133 ? 5'h7 : _T_719; // @[Lookup.scala 33:37]
  wire [4:0] _T_721 = _T_131 ? 5'h6 : _T_720; // @[Lookup.scala 33:37]
  wire [4:0] rvcImmType = _T_129 ? 5'he : _T_721; // @[Lookup.scala 33:37]
  wire [3:0] _T_722 = _T_193 ? 4'h9 : 4'h0; // @[Lookup.scala 33:37]
  wire [3:0] _T_723 = _T_191 ? 4'h9 : _T_722; // @[Lookup.scala 33:37]
  wire [3:0] _T_724 = _T_189 ? 4'h2 : _T_723; // @[Lookup.scala 33:37]
  wire [3:0] _T_725 = _T_187 ? 4'h4 : _T_724; // @[Lookup.scala 33:37]
  wire [3:0] _T_726 = _T_185 ? 4'h0 : _T_725; // @[Lookup.scala 33:37]
  wire [3:0] _T_727 = _T_183 ? 4'h5 : _T_726; // @[Lookup.scala 33:37]
  wire [3:0] _T_728 = _T_181 ? 4'h4 : _T_727; // @[Lookup.scala 33:37]
  wire [3:0] _T_729 = _T_179 ? 4'h9 : _T_728; // @[Lookup.scala 33:37]
  wire [3:0] _T_730 = _T_177 ? 4'h9 : _T_729; // @[Lookup.scala 33:37]
  wire [3:0] _T_731 = _T_175 ? 4'h2 : _T_730; // @[Lookup.scala 33:37]
  wire [3:0] _T_732 = _T_173 ? 4'h6 : _T_731; // @[Lookup.scala 33:37]
  wire [3:0] _T_733 = _T_171 ? 4'h6 : _T_732; // @[Lookup.scala 33:37]
  wire [3:0] _T_734 = _T_169 ? 4'h0 : _T_733; // @[Lookup.scala 33:37]
  wire [3:0] _T_735 = _T_167 ? 4'h6 : _T_734; // @[Lookup.scala 33:37]
  wire [3:0] _T_736 = _T_165 ? 4'h6 : _T_735; // @[Lookup.scala 33:37]
  wire [3:0] _T_737 = _T_163 ? 4'h6 : _T_736; // @[Lookup.scala 33:37]
  wire [3:0] _T_738 = _T_161 ? 4'h6 : _T_737; // @[Lookup.scala 33:37]
  wire [3:0] _T_739 = _T_159 ? 4'h6 : _T_738; // @[Lookup.scala 33:37]
  wire [3:0] _T_740 = _T_157 ? 4'h6 : _T_739; // @[Lookup.scala 33:37]
  wire [3:0] _T_741 = _T_155 ? 4'h6 : _T_740; // @[Lookup.scala 33:37]
  wire [3:0] _T_742 = _T_153 ? 4'h6 : _T_741; // @[Lookup.scala 33:37]
  wire [3:0] _T_743 = _T_151 ? 4'h6 : _T_742; // @[Lookup.scala 33:37]
  wire [3:0] _T_744 = _T_149 ? 4'h0 : _T_743; // @[Lookup.scala 33:37]
  wire [3:0] _T_745 = _T_147 ? 4'h9 : _T_744; // @[Lookup.scala 33:37]
  wire [3:0] _T_746 = _T_145 ? 4'h0 : _T_745; // @[Lookup.scala 33:37]
  wire [3:0] _T_747 = _T_143 ? 4'h2 : _T_746; // @[Lookup.scala 33:37]
  wire [3:0] _T_748 = _T_141 ? 4'h2 : _T_747; // @[Lookup.scala 33:37]
  wire [3:0] _T_749 = _T_139 ? 4'h0 : _T_748; // @[Lookup.scala 33:37]
  wire [3:0] _T_750 = _T_137 ? 4'h6 : _T_749; // @[Lookup.scala 33:37]
  wire [3:0] _T_751 = _T_135 ? 4'h6 : _T_750; // @[Lookup.scala 33:37]
  wire [3:0] _T_752 = _T_133 ? 4'h6 : _T_751; // @[Lookup.scala 33:37]
  wire [3:0] _T_753 = _T_131 ? 4'h6 : _T_752; // @[Lookup.scala 33:37]
  wire [3:0] rvcSrc1Type = _T_129 ? 4'h9 : _T_753; // @[Lookup.scala 33:37]
  wire [2:0] _T_754 = _T_193 ? 3'h5 : 3'h0; // @[Lookup.scala 33:37]
  wire [2:0] _T_755 = _T_191 ? 3'h5 : _T_754; // @[Lookup.scala 33:37]
  wire [2:0] _T_756 = _T_189 ? 3'h5 : _T_755; // @[Lookup.scala 33:37]
  wire [2:0] _T_757 = _T_187 ? 3'h0 : _T_756; // @[Lookup.scala 33:37]
  wire [2:0] _T_758 = _T_185 ? 3'h0 : _T_757; // @[Lookup.scala 33:37]
  wire [2:0] _T_759 = _T_183 ? 3'h0 : _T_758; // @[Lookup.scala 33:37]
  wire [2:0] _T_760 = _T_181 ? 3'h0 : _T_759; // @[Lookup.scala 33:37]
  wire [2:0] _T_761 = _T_179 ? 3'h0 : _T_760; // @[Lookup.scala 33:37]
  wire [2:0] _T_762 = _T_177 ? 3'h0 : _T_761; // @[Lookup.scala 33:37]
  wire [2:0] _T_763 = _T_175 ? 3'h0 : _T_762; // @[Lookup.scala 33:37]
  wire [2:0] _T_764 = _T_173 ? 3'h0 : _T_763; // @[Lookup.scala 33:37]
  wire [2:0] _T_765 = _T_171 ? 3'h0 : _T_764; // @[Lookup.scala 33:37]
  wire [2:0] _T_766 = _T_169 ? 3'h0 : _T_765; // @[Lookup.scala 33:37]
  wire [2:0] _T_767 = _T_167 ? 3'h7 : _T_766; // @[Lookup.scala 33:37]
  wire [2:0] _T_768 = _T_165 ? 3'h7 : _T_767; // @[Lookup.scala 33:37]
  wire [2:0] _T_769 = _T_163 ? 3'h7 : _T_768; // @[Lookup.scala 33:37]
  wire [2:0] _T_770 = _T_161 ? 3'h7 : _T_769; // @[Lookup.scala 33:37]
  wire [2:0] _T_771 = _T_159 ? 3'h7 : _T_770; // @[Lookup.scala 33:37]
  wire [2:0] _T_772 = _T_157 ? 3'h7 : _T_771; // @[Lookup.scala 33:37]
  wire [2:0] _T_773 = _T_155 ? 3'h0 : _T_772; // @[Lookup.scala 33:37]
  wire [2:0] _T_774 = _T_153 ? 3'h0 : _T_773; // @[Lookup.scala 33:37]
  wire [2:0] _T_775 = _T_151 ? 3'h0 : _T_774; // @[Lookup.scala 33:37]
  wire [2:0] _T_776 = _T_149 ? 3'h0 : _T_775; // @[Lookup.scala 33:37]
  wire [2:0] _T_777 = _T_147 ? 3'h0 : _T_776; // @[Lookup.scala 33:37]
  wire [2:0] _T_778 = _T_145 ? 3'h0 : _T_777; // @[Lookup.scala 33:37]
  wire [2:0] _T_779 = _T_143 ? 3'h0 : _T_778; // @[Lookup.scala 33:37]
  wire [2:0] _T_780 = _T_141 ? 3'h0 : _T_779; // @[Lookup.scala 33:37]
  wire [2:0] _T_781 = _T_139 ? 3'h0 : _T_780; // @[Lookup.scala 33:37]
  wire [2:0] _T_782 = _T_137 ? 3'h7 : _T_781; // @[Lookup.scala 33:37]
  wire [2:0] _T_783 = _T_135 ? 3'h7 : _T_782; // @[Lookup.scala 33:37]
  wire [2:0] _T_784 = _T_133 ? 3'h0 : _T_783; // @[Lookup.scala 33:37]
  wire [2:0] _T_785 = _T_131 ? 3'h0 : _T_784; // @[Lookup.scala 33:37]
  wire [2:0] rvcSrc2Type = _T_129 ? 3'h0 : _T_785; // @[Lookup.scala 33:37]
  wire [1:0] _T_788 = _T_189 ? 2'h2 : 2'h0; // @[Lookup.scala 33:37]
  wire [3:0] _T_789 = _T_187 ? 4'h8 : {{2'd0}, _T_788}; // @[Lookup.scala 33:37]
  wire [3:0] _T_790 = _T_185 ? 4'h0 : _T_789; // @[Lookup.scala 33:37]
  wire [3:0] _T_791 = _T_183 ? 4'h2 : _T_790; // @[Lookup.scala 33:37]
  wire [3:0] _T_792 = _T_181 ? 4'h0 : _T_791; // @[Lookup.scala 33:37]
  wire [3:0] _T_793 = _T_179 ? 4'h2 : _T_792; // @[Lookup.scala 33:37]
  wire [3:0] _T_794 = _T_177 ? 4'h2 : _T_793; // @[Lookup.scala 33:37]
  wire [3:0] _T_795 = _T_175 ? 4'h2 : _T_794; // @[Lookup.scala 33:37]
  wire [3:0] _T_796 = _T_173 ? 4'h0 : _T_795; // @[Lookup.scala 33:37]
  wire [3:0] _T_797 = _T_171 ? 4'h0 : _T_796; // @[Lookup.scala 33:37]
  wire [3:0] _T_798 = _T_169 ? 4'h0 : _T_797; // @[Lookup.scala 33:37]
  wire [3:0] _T_799 = _T_167 ? 4'h6 : _T_798; // @[Lookup.scala 33:37]
  wire [3:0] _T_800 = _T_165 ? 4'h6 : _T_799; // @[Lookup.scala 33:37]
  wire [3:0] _T_801 = _T_163 ? 4'h6 : _T_800; // @[Lookup.scala 33:37]
  wire [3:0] _T_802 = _T_161 ? 4'h6 : _T_801; // @[Lookup.scala 33:37]
  wire [3:0] _T_803 = _T_159 ? 4'h6 : _T_802; // @[Lookup.scala 33:37]
  wire [3:0] _T_804 = _T_157 ? 4'h6 : _T_803; // @[Lookup.scala 33:37]
  wire [3:0] _T_805 = _T_155 ? 4'h6 : _T_804; // @[Lookup.scala 33:37]
  wire [3:0] _T_806 = _T_153 ? 4'h6 : _T_805; // @[Lookup.scala 33:37]
  wire [3:0] _T_807 = _T_151 ? 4'h6 : _T_806; // @[Lookup.scala 33:37]
  wire [3:0] _T_808 = _T_149 ? 4'h2 : _T_807; // @[Lookup.scala 33:37]
  wire [3:0] _T_809 = _T_147 ? 4'h9 : _T_808; // @[Lookup.scala 33:37]
  wire [3:0] _T_810 = _T_145 ? 4'h2 : _T_809; // @[Lookup.scala 33:37]
  wire [3:0] _T_811 = _T_143 ? 4'h2 : _T_810; // @[Lookup.scala 33:37]
  wire [3:0] _T_812 = _T_141 ? 4'h2 : _T_811; // @[Lookup.scala 33:37]
  wire [3:0] _T_813 = _T_139 ? 4'h0 : _T_812; // @[Lookup.scala 33:37]
  wire [3:0] _T_814 = _T_137 ? 4'h0 : _T_813; // @[Lookup.scala 33:37]
  wire [3:0] _T_815 = _T_135 ? 4'h0 : _T_814; // @[Lookup.scala 33:37]
  wire [3:0] _T_816 = _T_133 ? 4'h7 : _T_815; // @[Lookup.scala 33:37]
  wire [3:0] _T_817 = _T_131 ? 4'h7 : _T_816; // @[Lookup.scala 33:37]
  wire [3:0] rvcDestType = _T_129 ? 4'h7 : _T_817; // @[Lookup.scala 33:37]
  wire  _T_818 = 4'h4 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_820 = 4'h2 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_821 = 4'hf == instrType; // @[LookupTree.scala 24:34]
  wire  _T_822 = 4'h1 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_823 = 4'h6 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_824 = 4'h7 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_825 = 4'h0 == instrType; // @[LookupTree.scala 24:34]
  wire  _T_839 = _T_823 | _T_824; // @[Mux.scala 27:72]
  wire  src1Type = _T_839 | _T_825; // @[Mux.scala 27:72]
  wire  _T_861 = _T_818 | _T_823; // @[Mux.scala 27:72]
  wire  _T_862 = _T_861 | _T_824; // @[Mux.scala 27:72]
  wire  src2Type = _T_862 | _T_825; // @[Mux.scala 27:72]
  wire [4:0] rs = io_in_bits_instr[19:15]; // @[IDU.scala 60:28]
  wire [4:0] rt = io_in_bits_instr[24:20]; // @[IDU.scala 60:43]
  wire [4:0] rd = io_in_bits_instr[11:7]; // @[IDU.scala 60:58]
  wire [4:0] rs2 = io_in_bits_instr[6:2]; // @[IDU.scala 63:24]
  wire  _T_865 = 3'h0 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_866 = 3'h1 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_867 = 3'h2 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_868 = 3'h3 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_869 = 3'h4 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_870 = 3'h5 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_871 = 3'h6 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire  _T_872 = 3'h7 == io_in_bits_instr[9:7]; // @[LookupTree.scala 24:34]
  wire [3:0] _T_873 = _T_865 ? 4'h8 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_874 = _T_866 ? 4'h9 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_875 = _T_867 ? 4'ha : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_876 = _T_868 ? 4'hb : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_877 = _T_869 ? 4'hc : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_878 = _T_870 ? 4'hd : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_879 = _T_871 ? 4'he : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_880 = _T_872 ? 4'hf : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_881 = _T_873 | _T_874; // @[Mux.scala 27:72]
  wire [3:0] _T_882 = _T_881 | _T_875; // @[Mux.scala 27:72]
  wire [3:0] _T_883 = _T_882 | _T_876; // @[Mux.scala 27:72]
  wire [3:0] _T_884 = _T_883 | _T_877; // @[Mux.scala 27:72]
  wire [3:0] _T_885 = _T_884 | _T_878; // @[Mux.scala 27:72]
  wire [3:0] _T_886 = _T_885 | _T_879; // @[Mux.scala 27:72]
  wire [3:0] rs1p = _T_886 | _T_880; // @[Mux.scala 27:72]
  wire  _T_889 = 3'h0 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_890 = 3'h1 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_891 = 3'h2 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_892 = 3'h3 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_893 = 3'h4 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_894 = 3'h5 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_895 = 3'h6 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire  _T_896 = 3'h7 == io_in_bits_instr[4:2]; // @[LookupTree.scala 24:34]
  wire [3:0] _T_897 = _T_889 ? 4'h8 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_898 = _T_890 ? 4'h9 : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_899 = _T_891 ? 4'ha : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_900 = _T_892 ? 4'hb : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_901 = _T_893 ? 4'hc : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_902 = _T_894 ? 4'hd : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_903 = _T_895 ? 4'he : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_904 = _T_896 ? 4'hf : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_905 = _T_897 | _T_898; // @[Mux.scala 27:72]
  wire [3:0] _T_906 = _T_905 | _T_899; // @[Mux.scala 27:72]
  wire [3:0] _T_907 = _T_906 | _T_900; // @[Mux.scala 27:72]
  wire [3:0] _T_908 = _T_907 | _T_901; // @[Mux.scala 27:72]
  wire [3:0] _T_909 = _T_908 | _T_902; // @[Mux.scala 27:72]
  wire [3:0] _T_910 = _T_909 | _T_903; // @[Mux.scala 27:72]
  wire [3:0] rs2p = _T_910 | _T_904; // @[Mux.scala 27:72]
  wire [5:0] rvc_shamt = {io_in_bits_instr[12],rs2}; // @[Cat.scala 29:58]
  wire  _T_915 = 4'h3 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_916 = 4'h1 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_917 = 4'h2 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_918 = 4'h4 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_919 = 4'h5 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_920 = 4'h6 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_921 = 4'h7 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_922 = 4'h8 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire  _T_923 = 4'h9 == rvcSrc1Type; // @[LookupTree.scala 24:34]
  wire [4:0] _T_925 = _T_915 ? rs : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_926 = _T_916 ? rt : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_927 = _T_917 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_928 = _T_918 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_929 = _T_919 ? rs2 : 5'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_930 = _T_920 ? rs1p : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_931 = _T_921 ? rs2p : 4'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_933 = _T_923 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_935 = _T_925 | _T_926; // @[Mux.scala 27:72]
  wire [4:0] _T_936 = _T_935 | _T_927; // @[Mux.scala 27:72]
  wire [4:0] _T_937 = _T_936 | _T_928; // @[Mux.scala 27:72]
  wire [4:0] _T_938 = _T_937 | _T_929; // @[Mux.scala 27:72]
  wire [4:0] _GEN_5 = {{1'd0}, _T_930}; // @[Mux.scala 27:72]
  wire [4:0] _T_939 = _T_938 | _GEN_5; // @[Mux.scala 27:72]
  wire [4:0] _GEN_6 = {{1'd0}, _T_931}; // @[Mux.scala 27:72]
  wire [4:0] _T_940 = _T_939 | _GEN_6; // @[Mux.scala 27:72]
  wire [4:0] _GEN_7 = {{4'd0}, _T_922}; // @[Mux.scala 27:72]
  wire [4:0] _T_941 = _T_940 | _GEN_7; // @[Mux.scala 27:72]
  wire [4:0] _GEN_8 = {{3'd0}, _T_933}; // @[Mux.scala 27:72]
  wire [4:0] rvc_src1 = _T_941 | _GEN_8; // @[Mux.scala 27:72]
  wire  _T_944 = 3'h3 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_945 = 3'h1 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_946 = 3'h2 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_947 = 3'h4 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_948 = 3'h5 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_949 = 3'h6 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire  _T_950 = 3'h7 == rvcSrc2Type; // @[LookupTree.scala 24:34]
  wire [3:0] _GEN_9 = {{1'd0}, rvcSrc2Type}; // @[LookupTree.scala 24:34]
  wire  _T_951 = 4'h8 == _GEN_9; // @[LookupTree.scala 24:34]
  wire  _T_952 = 4'h9 == _GEN_9; // @[LookupTree.scala 24:34]
  wire [4:0] _T_954 = _T_944 ? rs : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_955 = _T_945 ? rt : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_956 = _T_946 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_957 = _T_947 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_958 = _T_948 ? rs2 : 5'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_959 = _T_949 ? rs1p : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_960 = _T_950 ? rs2p : 4'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_962 = _T_952 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_964 = _T_954 | _T_955; // @[Mux.scala 27:72]
  wire [4:0] _T_965 = _T_964 | _T_956; // @[Mux.scala 27:72]
  wire [4:0] _T_966 = _T_965 | _T_957; // @[Mux.scala 27:72]
  wire [4:0] _T_967 = _T_966 | _T_958; // @[Mux.scala 27:72]
  wire [4:0] _GEN_11 = {{1'd0}, _T_959}; // @[Mux.scala 27:72]
  wire [4:0] _T_968 = _T_967 | _GEN_11; // @[Mux.scala 27:72]
  wire [4:0] _GEN_12 = {{1'd0}, _T_960}; // @[Mux.scala 27:72]
  wire [4:0] _T_969 = _T_968 | _GEN_12; // @[Mux.scala 27:72]
  wire [4:0] _GEN_13 = {{4'd0}, _T_951}; // @[Mux.scala 27:72]
  wire [4:0] _T_970 = _T_969 | _GEN_13; // @[Mux.scala 27:72]
  wire [4:0] _GEN_14 = {{3'd0}, _T_962}; // @[Mux.scala 27:72]
  wire [4:0] rvc_src2 = _T_970 | _GEN_14; // @[Mux.scala 27:72]
  wire  _T_973 = 4'h3 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_974 = 4'h1 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_975 = 4'h2 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_976 = 4'h4 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_977 = 4'h5 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_978 = 4'h6 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_979 = 4'h7 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_980 = 4'h8 == rvcDestType; // @[LookupTree.scala 24:34]
  wire  _T_981 = 4'h9 == rvcDestType; // @[LookupTree.scala 24:34]
  wire [4:0] _T_983 = _T_973 ? rs : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_984 = _T_974 ? rt : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_985 = _T_975 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_986 = _T_976 ? rd : 5'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_987 = _T_977 ? rs2 : 5'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_988 = _T_978 ? rs1p : 4'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_989 = _T_979 ? rs2p : 4'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_991 = _T_981 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [4:0] _T_993 = _T_983 | _T_984; // @[Mux.scala 27:72]
  wire [4:0] _T_994 = _T_993 | _T_985; // @[Mux.scala 27:72]
  wire [4:0] _T_995 = _T_994 | _T_986; // @[Mux.scala 27:72]
  wire [4:0] _T_996 = _T_995 | _T_987; // @[Mux.scala 27:72]
  wire [4:0] _GEN_15 = {{1'd0}, _T_988}; // @[Mux.scala 27:72]
  wire [4:0] _T_997 = _T_996 | _GEN_15; // @[Mux.scala 27:72]
  wire [4:0] _GEN_16 = {{1'd0}, _T_989}; // @[Mux.scala 27:72]
  wire [4:0] _T_998 = _T_997 | _GEN_16; // @[Mux.scala 27:72]
  wire [4:0] _GEN_17 = {{4'd0}, _T_980}; // @[Mux.scala 27:72]
  wire [4:0] _T_999 = _T_998 | _GEN_17; // @[Mux.scala 27:72]
  wire [4:0] _GEN_18 = {{3'd0}, _T_991}; // @[Mux.scala 27:72]
  wire [4:0] rvc_dest = _T_999 | _GEN_18; // @[Mux.scala 27:72]
  wire [4:0] rfSrc1 = isRVC ? rvc_src1 : rs; // @[IDU.scala 87:19]
  wire [4:0] rfSrc2 = isRVC ? rvc_src2 : rt; // @[IDU.scala 88:19]
  wire [4:0] rfDest = isRVC ? rvc_dest : rd; // @[IDU.scala 89:19]
  wire  _T_1003 = ~src2Type; // @[IDU.scala 93:43]
  wire [51:0] _T_1011 = io_in_bits_instr[31] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1012 = {_T_1011,io_in_bits_instr[31:20]}; // @[Cat.scala 29:58]
  wire [11:0] _T_1015 = {io_in_bits_instr[31:25],rd}; // @[Cat.scala 29:58]
  wire [51:0] _T_1018 = _T_1015[11] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1019 = {_T_1018,io_in_bits_instr[31:25],rd}; // @[Cat.scala 29:58]
  wire [12:0] _T_1034 = {io_in_bits_instr[31],io_in_bits_instr[7],io_in_bits_instr[30:25],io_in_bits_instr[11:8],1'h0}; // @[Cat.scala 29:58]
  wire [50:0] _T_1037 = _T_1034[12] ? 51'h7ffffffffffff : 51'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1038 = {_T_1037,io_in_bits_instr[31],io_in_bits_instr[7],io_in_bits_instr[30:25],io_in_bits_instr[11:8],1'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_1040 = {io_in_bits_instr[31:12],12'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_1043 = _T_1040[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1044 = {_T_1043,io_in_bits_instr[31:12],12'h0}; // @[Cat.scala 29:58]
  wire [20:0] _T_1052 = {io_in_bits_instr[31],io_in_bits_instr[19:12],io_in_bits_instr[20],io_in_bits_instr[30:21],1'h0}; // @[Cat.scala 29:58]
  wire [42:0] _T_1055 = _T_1052[20] ? 43'h7ffffffffff : 43'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1056 = {_T_1055,io_in_bits_instr[31],io_in_bits_instr[19:12],io_in_bits_instr[20],io_in_bits_instr[30:21],1'h0}; // @[Cat.scala 29:58]
  wire [63:0] _T_1063 = _T_818 ? _T_1012 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1064 = _T_820 ? _T_1019 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1065 = _T_821 ? _T_1019 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1066 = _T_822 ? _T_1038 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1067 = _T_823 ? _T_1044 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1068 = _T_824 ? _T_1056 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1069 = _T_1063 | _T_1064; // @[Mux.scala 27:72]
  wire [63:0] _T_1070 = _T_1069 | _T_1065; // @[Mux.scala 27:72]
  wire [63:0] _T_1071 = _T_1070 | _T_1066; // @[Mux.scala 27:72]
  wire [63:0] _T_1072 = _T_1071 | _T_1067; // @[Mux.scala 27:72]
  wire [63:0] imm = _T_1072 | _T_1068; // @[Mux.scala 27:72]
  wire [63:0] _T_1080 = {56'h0,io_in_bits_instr[3:2],io_in_bits_instr[12],io_in_bits_instr[6:4],2'h0}; // @[Cat.scala 29:58]
  wire [63:0] _T_1087 = {55'h0,io_in_bits_instr[4:2],io_in_bits_instr[12],io_in_bits_instr[6:5],3'h0}; // @[Cat.scala 29:58]
  wire [63:0] _T_1092 = {56'h0,io_in_bits_instr[8:7],io_in_bits_instr[12:9],2'h0}; // @[Cat.scala 29:58]
  wire [63:0] _T_1097 = {55'h0,io_in_bits_instr[9:7],io_in_bits_instr[12:10],3'h0}; // @[Cat.scala 29:58]
  wire [63:0] _T_1104 = {57'h0,io_in_bits_instr[5],io_in_bits_instr[12:10],io_in_bits_instr[6],2'h0}; // @[Cat.scala 29:58]
  wire [63:0] _T_1109 = {56'h0,io_in_bits_instr[6:5],io_in_bits_instr[12:10],3'h0}; // @[Cat.scala 29:58]
  wire [11:0] _T_1137 = {io_in_bits_instr[12],io_in_bits_instr[8],io_in_bits_instr[10:9],io_in_bits_instr[6],io_in_bits_instr[7],io_in_bits_instr[2],io_in_bits_instr[11],io_in_bits_instr[5:3],1'h0}; // @[Cat.scala 29:58]
  wire [51:0] _T_1140 = _T_1137[11] ? 52'hfffffffffffff : 52'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1141 = {_T_1140,io_in_bits_instr[12],io_in_bits_instr[8],io_in_bits_instr[10:9],io_in_bits_instr[6],io_in_bits_instr[7],io_in_bits_instr[2],io_in_bits_instr[11],io_in_bits_instr[5:3],1'h0}; // @[Cat.scala 29:58]
  wire [8:0] _T_1151 = {io_in_bits_instr[12],io_in_bits_instr[6:5],io_in_bits_instr[2],io_in_bits_instr[11:10],io_in_bits_instr[4:3],1'h0}; // @[Cat.scala 29:58]
  wire [54:0] _T_1154 = _T_1151[8] ? 55'h7fffffffffffff : 55'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1155 = {_T_1154,io_in_bits_instr[12],io_in_bits_instr[6:5],io_in_bits_instr[2],io_in_bits_instr[11:10],io_in_bits_instr[4:3],1'h0}; // @[Cat.scala 29:58]
  wire [57:0] _T_1161 = rvc_shamt[5] ? 58'h3ffffffffffffff : 58'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1162 = {_T_1161,io_in_bits_instr[12],rs2}; // @[Cat.scala 29:58]
  wire [17:0] _T_1166 = {io_in_bits_instr[12],rs2,12'h0}; // @[Cat.scala 29:58]
  wire [45:0] _T_1169 = _T_1166[17] ? 46'h3fffffffffff : 46'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1170 = {_T_1169,io_in_bits_instr[12],rs2,12'h0}; // @[Cat.scala 29:58]
  wire [9:0] _T_1187 = {io_in_bits_instr[12],io_in_bits_instr[4:3],io_in_bits_instr[5],io_in_bits_instr[2],io_in_bits_instr[6],4'h0}; // @[Cat.scala 29:58]
  wire [53:0] _T_1190 = _T_1187[9] ? 54'h3fffffffffffff : 54'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_1191 = {_T_1190,io_in_bits_instr[12],io_in_bits_instr[4:3],io_in_bits_instr[5],io_in_bits_instr[2],io_in_bits_instr[6],4'h0}; // @[Cat.scala 29:58]
  wire [63:0] _T_1200 = {54'h0,io_in_bits_instr[10:7],io_in_bits_instr[12:11],io_in_bits_instr[5],io_in_bits_instr[6],2'h0}; // @[Cat.scala 29:58]
  wire  _T_1202 = 5'h0 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1203 = 5'h1 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1204 = 5'h2 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1205 = 5'h3 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1206 = 5'h4 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1207 = 5'h5 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1208 = 5'h6 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1209 = 5'h7 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1210 = 5'h8 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1211 = 5'h9 == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1212 = 5'ha == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1213 = 5'hb == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1214 = 5'hc == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1215 = 5'hd == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1216 = 5'he == rvcImmType; // @[LookupTree.scala 24:34]
  wire  _T_1217 = 5'hf == rvcImmType; // @[LookupTree.scala 24:34]
  wire [63:0] _T_1219 = _T_1202 ? _T_1080 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1220 = _T_1203 ? _T_1087 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1221 = _T_1204 ? _T_1092 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1222 = _T_1205 ? _T_1097 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1223 = _T_1206 ? _T_1104 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1224 = _T_1207 ? _T_1109 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1225 = _T_1208 ? _T_1104 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1226 = _T_1209 ? _T_1109 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1227 = _T_1210 ? _T_1141 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1228 = _T_1211 ? _T_1155 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1229 = _T_1212 ? _T_1162 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1230 = _T_1213 ? _T_1170 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1231 = _T_1214 ? _T_1162 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1232 = _T_1215 ? _T_1191 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1233 = _T_1216 ? _T_1200 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1234 = _T_1217 ? 64'h1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_1236 = _T_1219 | _T_1220; // @[Mux.scala 27:72]
  wire [63:0] _T_1237 = _T_1236 | _T_1221; // @[Mux.scala 27:72]
  wire [63:0] _T_1238 = _T_1237 | _T_1222; // @[Mux.scala 27:72]
  wire [63:0] _T_1239 = _T_1238 | _T_1223; // @[Mux.scala 27:72]
  wire [63:0] _T_1240 = _T_1239 | _T_1224; // @[Mux.scala 27:72]
  wire [63:0] _T_1241 = _T_1240 | _T_1225; // @[Mux.scala 27:72]
  wire [63:0] _T_1242 = _T_1241 | _T_1226; // @[Mux.scala 27:72]
  wire [63:0] _T_1243 = _T_1242 | _T_1227; // @[Mux.scala 27:72]
  wire [63:0] _T_1244 = _T_1243 | _T_1228; // @[Mux.scala 27:72]
  wire [63:0] _T_1245 = _T_1244 | _T_1229; // @[Mux.scala 27:72]
  wire [63:0] _T_1246 = _T_1245 | _T_1230; // @[Mux.scala 27:72]
  wire [63:0] _T_1247 = _T_1246 | _T_1231; // @[Mux.scala 27:72]
  wire [63:0] _T_1248 = _T_1247 | _T_1232; // @[Mux.scala 27:72]
  wire [63:0] _T_1249 = _T_1248 | _T_1233; // @[Mux.scala 27:72]
  wire [63:0] immrvc = _T_1249 | _T_1234; // @[Mux.scala 27:72]
  wire  _T_1252 = fuType == 3'h0; // @[IDU.scala 130:16]
  wire  _T_1253 = rfDest == 5'h1; // @[IDU.scala 131:34]
  wire  _T_1254 = rfDest == 5'h5; // @[IDU.scala 131:49]
  wire  _T_1255 = _T_1253 | _T_1254; // @[IDU.scala 131:42]
  wire  _T_1256 = fuOpType == 7'h58; // @[IDU.scala 132:38]
  wire  _T_1257 = _T_1255 & _T_1256; // @[IDU.scala 132:26]
  wire [6:0] _GEN_0 = _T_1257 ? 7'h5c : fuOpType; // @[IDU.scala 132:57]
  wire  _T_1258 = fuOpType == 7'h5a; // @[IDU.scala 133:20]
  wire  _T_1259 = rfSrc1 == 5'h1; // @[IDU.scala 131:34]
  wire  _T_1260 = rfSrc1 == 5'h5; // @[IDU.scala 131:49]
  wire  _T_1261 = _T_1259 | _T_1260; // @[IDU.scala 131:42]
  wire [6:0] _GEN_1 = _T_1261 ? 7'h5e : _GEN_0; // @[IDU.scala 134:29]
  wire [6:0] _GEN_2 = _T_1255 ? 7'h5c : _GEN_1; // @[IDU.scala 135:29]
  wire [6:0] _GEN_3 = _T_1258 ? _GEN_2 : _GEN_0; // @[IDU.scala 133:40]
  wire  _T_1266 = io_in_bits_instr[6:0] == 7'h37; // @[IDU.scala 139:47]
  wire  _T_1278 = ~io_in_valid; // @[IDU.scala 160:18]
  wire  _T_1279 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_1280 = ~hasIntr; // @[IDU.scala 160:51]
  wire  _T_1281 = _T_1279 & _T_1280; // @[IDU.scala 160:48]
  wire  _T_1306 = instrType == 4'h0; // @[IDU.scala 176:59]
  wire  _T_1308 = _T_1306 & _T_1280; // @[IDU.scala 176:70]
  wire  _T_1311 = |io_in_bits_pc[38:32]; // @[IDU.scala 179:94]
  wire  _T_1312 = ~DTLBENABLE; // @[IDU.scala 179:101]
  assign io_in_ready = _T_1278 | _T_1281; // @[IDU.scala 160:15]
  assign io_out_valid = io_in_valid; // @[IDU.scala 159:16]
  assign io_out_bits_cf_instr = io_in_bits_instr; // @[IDU.scala 161:18]
  assign io_out_bits_cf_pc = io_in_bits_pc; // @[IDU.scala 161:18]
  assign io_out_bits_cf_pnpc = io_in_bits_pnpc; // @[IDU.scala 161:18]
  assign io_out_bits_cf_exceptionVec_1 = _T_1311 & _T_1312; // @[IDU.scala 161:18 IDU.scala 175:37 IDU.scala 179:51]
  assign io_out_bits_cf_exceptionVec_2 = _T_1308 & io_in_valid; // @[IDU.scala 161:18 IDU.scala 175:37 IDU.scala 176:45]
  assign io_out_bits_cf_exceptionVec_12 = io_in_bits_exceptionVec_12; // @[IDU.scala 161:18 IDU.scala 175:37 IDU.scala 177:47]
  assign io_out_bits_cf_intrVec_0 = intrVecIDU[0]; // @[IDU.scala 161:18 IDU.scala 169:68]
  assign io_out_bits_cf_intrVec_1 = intrVecIDU[1]; // @[IDU.scala 161:18 IDU.scala 169:68]
  assign io_out_bits_cf_intrVec_2 = intrVecIDU[2]; // @[IDU.scala 161:18 IDU.scala 169:68]
  assign io_out_bits_cf_intrVec_3 = intrVecIDU[3]; // @[IDU.scala 161:18 IDU.scala 169:68]
  assign io_out_bits_cf_intrVec_4 = intrVecIDU[4]; // @[IDU.scala 161:18 IDU.scala 169:68]
  assign io_out_bits_cf_intrVec_5 = intrVecIDU[5]; // @[IDU.scala 161:18 IDU.scala 169:68]
  assign io_out_bits_cf_intrVec_6 = intrVecIDU[6]; // @[IDU.scala 161:18 IDU.scala 169:68]
  assign io_out_bits_cf_intrVec_7 = intrVecIDU[7]; // @[IDU.scala 161:18 IDU.scala 169:68]
  assign io_out_bits_cf_intrVec_8 = intrVecIDU[8]; // @[IDU.scala 161:18 IDU.scala 169:68]
  assign io_out_bits_cf_intrVec_9 = intrVecIDU[9]; // @[IDU.scala 161:18 IDU.scala 169:68]
  assign io_out_bits_cf_intrVec_10 = intrVecIDU[10]; // @[IDU.scala 161:18 IDU.scala 169:68]
  assign io_out_bits_cf_intrVec_11 = intrVecIDU[11]; // @[IDU.scala 161:18 IDU.scala 169:68]
  assign io_out_bits_cf_brIdx = io_in_bits_brIdx; // @[IDU.scala 161:18]
  assign io_out_bits_cf_crossPageIPFFix = io_in_bits_crossPageIPFFix; // @[IDU.scala 161:18]
  assign io_out_bits_ctrl_src1Type = _T_1266 ? 1'h0 : src1Type; // @[IDU.scala 139:29]
  assign io_out_bits_ctrl_src2Type = _T_862 | _T_825; // @[IDU.scala 140:29]
  assign io_out_bits_ctrl_fuType = _T_618 ? 3'h3 : decodeList_1; // @[IDU.scala 44:27]
  assign io_out_bits_ctrl_fuOpType = _T_1252 ? _GEN_3 : fuOpType; // @[IDU.scala 45:29 IDU.scala 132:85 IDU.scala 134:57 IDU.scala 135:57]
  assign io_out_bits_ctrl_rfSrc1 = src1Type ? 5'h0 : rfSrc1; // @[IDU.scala 92:27]
  assign io_out_bits_ctrl_rfSrc2 = _T_1003 ? rfSrc2 : 5'h0; // @[IDU.scala 93:27]
  assign io_out_bits_ctrl_rfWen = instrType[2]; // @[IDU.scala 94:27]
  assign io_out_bits_ctrl_rfDest = instrType[2] ? rfDest : 5'h0; // @[IDU.scala 95:27]
  assign io_out_bits_data_imm = isRVC ? immrvc : imm; // @[IDU.scala 128:25]
endmodule
module Decoder_1(
  output        io_out_bits_cf_intrVec_0,
  output        io_out_bits_cf_intrVec_1,
  output        io_out_bits_cf_intrVec_2,
  output        io_out_bits_cf_intrVec_3,
  output        io_out_bits_cf_intrVec_4,
  output        io_out_bits_cf_intrVec_5,
  output        io_out_bits_cf_intrVec_6,
  output        io_out_bits_cf_intrVec_7,
  output        io_out_bits_cf_intrVec_8,
  output        io_out_bits_cf_intrVec_9,
  output        io_out_bits_cf_intrVec_10,
  output        io_out_bits_cf_intrVec_11,
  input  [11:0] intrVecIDU
);
  assign io_out_bits_cf_intrVec_0 = intrVecIDU[0]; // @[IDU.scala 161:18 IDU.scala 169:68]
  assign io_out_bits_cf_intrVec_1 = intrVecIDU[1]; // @[IDU.scala 161:18 IDU.scala 169:68]
  assign io_out_bits_cf_intrVec_2 = intrVecIDU[2]; // @[IDU.scala 161:18 IDU.scala 169:68]
  assign io_out_bits_cf_intrVec_3 = intrVecIDU[3]; // @[IDU.scala 161:18 IDU.scala 169:68]
  assign io_out_bits_cf_intrVec_4 = intrVecIDU[4]; // @[IDU.scala 161:18 IDU.scala 169:68]
  assign io_out_bits_cf_intrVec_5 = intrVecIDU[5]; // @[IDU.scala 161:18 IDU.scala 169:68]
  assign io_out_bits_cf_intrVec_6 = intrVecIDU[6]; // @[IDU.scala 161:18 IDU.scala 169:68]
  assign io_out_bits_cf_intrVec_7 = intrVecIDU[7]; // @[IDU.scala 161:18 IDU.scala 169:68]
  assign io_out_bits_cf_intrVec_8 = intrVecIDU[8]; // @[IDU.scala 161:18 IDU.scala 169:68]
  assign io_out_bits_cf_intrVec_9 = intrVecIDU[9]; // @[IDU.scala 161:18 IDU.scala 169:68]
  assign io_out_bits_cf_intrVec_10 = intrVecIDU[10]; // @[IDU.scala 161:18 IDU.scala 169:68]
  assign io_out_bits_cf_intrVec_11 = intrVecIDU[11]; // @[IDU.scala 161:18 IDU.scala 169:68]
endmodule
module IDU(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [63:0] io_in_0_bits_instr,
  input  [38:0] io_in_0_bits_pc,
  input  [38:0] io_in_0_bits_pnpc,
  input         io_in_0_bits_exceptionVec_12,
  input  [3:0]  io_in_0_bits_brIdx,
  input         io_in_0_bits_crossPageIPFFix,
  input         io_out_0_ready,
  output        io_out_0_valid,
  output [63:0] io_out_0_bits_cf_instr,
  output [38:0] io_out_0_bits_cf_pc,
  output [38:0] io_out_0_bits_cf_pnpc,
  output        io_out_0_bits_cf_exceptionVec_1,
  output        io_out_0_bits_cf_exceptionVec_2,
  output        io_out_0_bits_cf_exceptionVec_12,
  output        io_out_0_bits_cf_intrVec_0,
  output        io_out_0_bits_cf_intrVec_1,
  output        io_out_0_bits_cf_intrVec_2,
  output        io_out_0_bits_cf_intrVec_3,
  output        io_out_0_bits_cf_intrVec_4,
  output        io_out_0_bits_cf_intrVec_5,
  output        io_out_0_bits_cf_intrVec_6,
  output        io_out_0_bits_cf_intrVec_7,
  output        io_out_0_bits_cf_intrVec_8,
  output        io_out_0_bits_cf_intrVec_9,
  output        io_out_0_bits_cf_intrVec_10,
  output        io_out_0_bits_cf_intrVec_11,
  output [3:0]  io_out_0_bits_cf_brIdx,
  output        io_out_0_bits_cf_crossPageIPFFix,
  output        io_out_0_bits_ctrl_src1Type,
  output        io_out_0_bits_ctrl_src2Type,
  output [2:0]  io_out_0_bits_ctrl_fuType,
  output [6:0]  io_out_0_bits_ctrl_fuOpType,
  output [4:0]  io_out_0_bits_ctrl_rfSrc1,
  output [4:0]  io_out_0_bits_ctrl_rfSrc2,
  output        io_out_0_bits_ctrl_rfWen,
  output [4:0]  io_out_0_bits_ctrl_rfDest,
  output [63:0] io_out_0_bits_data_imm,
  output        io_out_1_bits_cf_intrVec_0,
  output        io_out_1_bits_cf_intrVec_1,
  output        io_out_1_bits_cf_intrVec_2,
  output        io_out_1_bits_cf_intrVec_3,
  output        io_out_1_bits_cf_intrVec_4,
  output        io_out_1_bits_cf_intrVec_5,
  output        io_out_1_bits_cf_intrVec_6,
  output        io_out_1_bits_cf_intrVec_7,
  output        io_out_1_bits_cf_intrVec_8,
  output        io_out_1_bits_cf_intrVec_9,
  output        io_out_1_bits_cf_intrVec_10,
  output        io_out_1_bits_cf_intrVec_11,
  input         vmEnable,
  input  [11:0] intrVec
);
  wire  decoder1_io_in_ready; // @[IDU.scala 194:25]
  wire  decoder1_io_in_valid; // @[IDU.scala 194:25]
  wire [63:0] decoder1_io_in_bits_instr; // @[IDU.scala 194:25]
  wire [38:0] decoder1_io_in_bits_pc; // @[IDU.scala 194:25]
  wire [38:0] decoder1_io_in_bits_pnpc; // @[IDU.scala 194:25]
  wire  decoder1_io_in_bits_exceptionVec_12; // @[IDU.scala 194:25]
  wire [3:0] decoder1_io_in_bits_brIdx; // @[IDU.scala 194:25]
  wire  decoder1_io_in_bits_crossPageIPFFix; // @[IDU.scala 194:25]
  wire  decoder1_io_out_ready; // @[IDU.scala 194:25]
  wire  decoder1_io_out_valid; // @[IDU.scala 194:25]
  wire [63:0] decoder1_io_out_bits_cf_instr; // @[IDU.scala 194:25]
  wire [38:0] decoder1_io_out_bits_cf_pc; // @[IDU.scala 194:25]
  wire [38:0] decoder1_io_out_bits_cf_pnpc; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_exceptionVec_1; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_exceptionVec_2; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_exceptionVec_12; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_intrVec_0; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_intrVec_1; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_intrVec_2; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_intrVec_3; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_intrVec_4; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_intrVec_5; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_intrVec_6; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_intrVec_7; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_intrVec_8; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_intrVec_9; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_intrVec_10; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_intrVec_11; // @[IDU.scala 194:25]
  wire [3:0] decoder1_io_out_bits_cf_brIdx; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_cf_crossPageIPFFix; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_ctrl_src1Type; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_ctrl_src2Type; // @[IDU.scala 194:25]
  wire [2:0] decoder1_io_out_bits_ctrl_fuType; // @[IDU.scala 194:25]
  wire [6:0] decoder1_io_out_bits_ctrl_fuOpType; // @[IDU.scala 194:25]
  wire [4:0] decoder1_io_out_bits_ctrl_rfSrc1; // @[IDU.scala 194:25]
  wire [4:0] decoder1_io_out_bits_ctrl_rfSrc2; // @[IDU.scala 194:25]
  wire  decoder1_io_out_bits_ctrl_rfWen; // @[IDU.scala 194:25]
  wire [4:0] decoder1_io_out_bits_ctrl_rfDest; // @[IDU.scala 194:25]
  wire [63:0] decoder1_io_out_bits_data_imm; // @[IDU.scala 194:25]
  wire  decoder1_DTLBENABLE; // @[IDU.scala 194:25]
  wire [11:0] decoder1_intrVecIDU; // @[IDU.scala 194:25]
  wire  decoder2_io_out_bits_cf_intrVec_0; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_cf_intrVec_1; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_cf_intrVec_2; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_cf_intrVec_3; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_cf_intrVec_4; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_cf_intrVec_5; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_cf_intrVec_6; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_cf_intrVec_7; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_cf_intrVec_8; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_cf_intrVec_9; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_cf_intrVec_10; // @[IDU.scala 195:25]
  wire  decoder2_io_out_bits_cf_intrVec_11; // @[IDU.scala 195:25]
  wire [11:0] decoder2_intrVecIDU; // @[IDU.scala 195:25]
  Decoder decoder1 ( // @[IDU.scala 194:25]
    .io_in_ready(decoder1_io_in_ready),
    .io_in_valid(decoder1_io_in_valid),
    .io_in_bits_instr(decoder1_io_in_bits_instr),
    .io_in_bits_pc(decoder1_io_in_bits_pc),
    .io_in_bits_pnpc(decoder1_io_in_bits_pnpc),
    .io_in_bits_exceptionVec_12(decoder1_io_in_bits_exceptionVec_12),
    .io_in_bits_brIdx(decoder1_io_in_bits_brIdx),
    .io_in_bits_crossPageIPFFix(decoder1_io_in_bits_crossPageIPFFix),
    .io_out_ready(decoder1_io_out_ready),
    .io_out_valid(decoder1_io_out_valid),
    .io_out_bits_cf_instr(decoder1_io_out_bits_cf_instr),
    .io_out_bits_cf_pc(decoder1_io_out_bits_cf_pc),
    .io_out_bits_cf_pnpc(decoder1_io_out_bits_cf_pnpc),
    .io_out_bits_cf_exceptionVec_1(decoder1_io_out_bits_cf_exceptionVec_1),
    .io_out_bits_cf_exceptionVec_2(decoder1_io_out_bits_cf_exceptionVec_2),
    .io_out_bits_cf_exceptionVec_12(decoder1_io_out_bits_cf_exceptionVec_12),
    .io_out_bits_cf_intrVec_0(decoder1_io_out_bits_cf_intrVec_0),
    .io_out_bits_cf_intrVec_1(decoder1_io_out_bits_cf_intrVec_1),
    .io_out_bits_cf_intrVec_2(decoder1_io_out_bits_cf_intrVec_2),
    .io_out_bits_cf_intrVec_3(decoder1_io_out_bits_cf_intrVec_3),
    .io_out_bits_cf_intrVec_4(decoder1_io_out_bits_cf_intrVec_4),
    .io_out_bits_cf_intrVec_5(decoder1_io_out_bits_cf_intrVec_5),
    .io_out_bits_cf_intrVec_6(decoder1_io_out_bits_cf_intrVec_6),
    .io_out_bits_cf_intrVec_7(decoder1_io_out_bits_cf_intrVec_7),
    .io_out_bits_cf_intrVec_8(decoder1_io_out_bits_cf_intrVec_8),
    .io_out_bits_cf_intrVec_9(decoder1_io_out_bits_cf_intrVec_9),
    .io_out_bits_cf_intrVec_10(decoder1_io_out_bits_cf_intrVec_10),
    .io_out_bits_cf_intrVec_11(decoder1_io_out_bits_cf_intrVec_11),
    .io_out_bits_cf_brIdx(decoder1_io_out_bits_cf_brIdx),
    .io_out_bits_cf_crossPageIPFFix(decoder1_io_out_bits_cf_crossPageIPFFix),
    .io_out_bits_ctrl_src1Type(decoder1_io_out_bits_ctrl_src1Type),
    .io_out_bits_ctrl_src2Type(decoder1_io_out_bits_ctrl_src2Type),
    .io_out_bits_ctrl_fuType(decoder1_io_out_bits_ctrl_fuType),
    .io_out_bits_ctrl_fuOpType(decoder1_io_out_bits_ctrl_fuOpType),
    .io_out_bits_ctrl_rfSrc1(decoder1_io_out_bits_ctrl_rfSrc1),
    .io_out_bits_ctrl_rfSrc2(decoder1_io_out_bits_ctrl_rfSrc2),
    .io_out_bits_ctrl_rfWen(decoder1_io_out_bits_ctrl_rfWen),
    .io_out_bits_ctrl_rfDest(decoder1_io_out_bits_ctrl_rfDest),
    .io_out_bits_data_imm(decoder1_io_out_bits_data_imm),
    .DTLBENABLE(decoder1_DTLBENABLE),
    .intrVecIDU(decoder1_intrVecIDU)
  );
  Decoder_1 decoder2 ( // @[IDU.scala 195:25]
    .io_out_bits_cf_intrVec_0(decoder2_io_out_bits_cf_intrVec_0),
    .io_out_bits_cf_intrVec_1(decoder2_io_out_bits_cf_intrVec_1),
    .io_out_bits_cf_intrVec_2(decoder2_io_out_bits_cf_intrVec_2),
    .io_out_bits_cf_intrVec_3(decoder2_io_out_bits_cf_intrVec_3),
    .io_out_bits_cf_intrVec_4(decoder2_io_out_bits_cf_intrVec_4),
    .io_out_bits_cf_intrVec_5(decoder2_io_out_bits_cf_intrVec_5),
    .io_out_bits_cf_intrVec_6(decoder2_io_out_bits_cf_intrVec_6),
    .io_out_bits_cf_intrVec_7(decoder2_io_out_bits_cf_intrVec_7),
    .io_out_bits_cf_intrVec_8(decoder2_io_out_bits_cf_intrVec_8),
    .io_out_bits_cf_intrVec_9(decoder2_io_out_bits_cf_intrVec_9),
    .io_out_bits_cf_intrVec_10(decoder2_io_out_bits_cf_intrVec_10),
    .io_out_bits_cf_intrVec_11(decoder2_io_out_bits_cf_intrVec_11),
    .intrVecIDU(decoder2_intrVecIDU)
  );
  assign io_in_0_ready = decoder1_io_in_ready; // @[IDU.scala 196:12]
  assign io_out_0_valid = decoder1_io_out_valid; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_instr = decoder1_io_out_bits_cf_instr; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_pc = decoder1_io_out_bits_cf_pc; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_pnpc = decoder1_io_out_bits_cf_pnpc; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_exceptionVec_1 = decoder1_io_out_bits_cf_exceptionVec_1; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_exceptionVec_2 = decoder1_io_out_bits_cf_exceptionVec_2; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_exceptionVec_12 = decoder1_io_out_bits_cf_exceptionVec_12; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_intrVec_0 = decoder1_io_out_bits_cf_intrVec_0; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_intrVec_1 = decoder1_io_out_bits_cf_intrVec_1; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_intrVec_2 = decoder1_io_out_bits_cf_intrVec_2; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_intrVec_3 = decoder1_io_out_bits_cf_intrVec_3; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_intrVec_4 = decoder1_io_out_bits_cf_intrVec_4; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_intrVec_5 = decoder1_io_out_bits_cf_intrVec_5; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_intrVec_6 = decoder1_io_out_bits_cf_intrVec_6; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_intrVec_7 = decoder1_io_out_bits_cf_intrVec_7; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_intrVec_8 = decoder1_io_out_bits_cf_intrVec_8; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_intrVec_9 = decoder1_io_out_bits_cf_intrVec_9; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_intrVec_10 = decoder1_io_out_bits_cf_intrVec_10; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_intrVec_11 = decoder1_io_out_bits_cf_intrVec_11; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_brIdx = decoder1_io_out_bits_cf_brIdx; // @[IDU.scala 198:13]
  assign io_out_0_bits_cf_crossPageIPFFix = decoder1_io_out_bits_cf_crossPageIPFFix; // @[IDU.scala 198:13]
  assign io_out_0_bits_ctrl_src1Type = decoder1_io_out_bits_ctrl_src1Type; // @[IDU.scala 198:13]
  assign io_out_0_bits_ctrl_src2Type = decoder1_io_out_bits_ctrl_src2Type; // @[IDU.scala 198:13]
  assign io_out_0_bits_ctrl_fuType = decoder1_io_out_bits_ctrl_fuType; // @[IDU.scala 198:13]
  assign io_out_0_bits_ctrl_fuOpType = decoder1_io_out_bits_ctrl_fuOpType; // @[IDU.scala 198:13]
  assign io_out_0_bits_ctrl_rfSrc1 = decoder1_io_out_bits_ctrl_rfSrc1; // @[IDU.scala 198:13]
  assign io_out_0_bits_ctrl_rfSrc2 = decoder1_io_out_bits_ctrl_rfSrc2; // @[IDU.scala 198:13]
  assign io_out_0_bits_ctrl_rfWen = decoder1_io_out_bits_ctrl_rfWen; // @[IDU.scala 198:13]
  assign io_out_0_bits_ctrl_rfDest = decoder1_io_out_bits_ctrl_rfDest; // @[IDU.scala 198:13]
  assign io_out_0_bits_data_imm = decoder1_io_out_bits_data_imm; // @[IDU.scala 198:13]
  assign io_out_1_bits_cf_intrVec_0 = decoder2_io_out_bits_cf_intrVec_0; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_intrVec_1 = decoder2_io_out_bits_cf_intrVec_1; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_intrVec_2 = decoder2_io_out_bits_cf_intrVec_2; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_intrVec_3 = decoder2_io_out_bits_cf_intrVec_3; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_intrVec_4 = decoder2_io_out_bits_cf_intrVec_4; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_intrVec_5 = decoder2_io_out_bits_cf_intrVec_5; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_intrVec_6 = decoder2_io_out_bits_cf_intrVec_6; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_intrVec_7 = decoder2_io_out_bits_cf_intrVec_7; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_intrVec_8 = decoder2_io_out_bits_cf_intrVec_8; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_intrVec_9 = decoder2_io_out_bits_cf_intrVec_9; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_intrVec_10 = decoder2_io_out_bits_cf_intrVec_10; // @[IDU.scala 199:13]
  assign io_out_1_bits_cf_intrVec_11 = decoder2_io_out_bits_cf_intrVec_11; // @[IDU.scala 199:13]
  assign decoder1_io_in_valid = io_in_0_valid; // @[IDU.scala 196:12]
  assign decoder1_io_in_bits_instr = io_in_0_bits_instr; // @[IDU.scala 196:12]
  assign decoder1_io_in_bits_pc = io_in_0_bits_pc; // @[IDU.scala 196:12]
  assign decoder1_io_in_bits_pnpc = io_in_0_bits_pnpc; // @[IDU.scala 196:12]
  assign decoder1_io_in_bits_exceptionVec_12 = io_in_0_bits_exceptionVec_12; // @[IDU.scala 196:12]
  assign decoder1_io_in_bits_brIdx = io_in_0_bits_brIdx; // @[IDU.scala 196:12]
  assign decoder1_io_in_bits_crossPageIPFFix = io_in_0_bits_crossPageIPFFix; // @[IDU.scala 196:12]
  assign decoder1_io_out_ready = io_out_0_ready; // @[IDU.scala 198:13]
  assign decoder1_DTLBENABLE = vmEnable;
  assign decoder1_intrVecIDU = intrVec;
  assign decoder2_intrVecIDU = intrVec;
endmodule
module FlushableQueue(
  input         clock,
  input         reset,
  output        io_enq_ready,
  input         io_enq_valid,
  input  [63:0] io_enq_bits_instr,
  input  [38:0] io_enq_bits_pc,
  input  [38:0] io_enq_bits_pnpc,
  input         io_enq_bits_exceptionVec_12,
  input  [3:0]  io_enq_bits_brIdx,
  input         io_deq_ready,
  output        io_deq_valid,
  output [63:0] io_deq_bits_instr,
  output [38:0] io_deq_bits_pc,
  output [38:0] io_deq_bits_pnpc,
  output        io_deq_bits_exceptionVec_12,
  output [3:0]  io_deq_bits_brIdx,
  input         io_flush
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] ram_instr [0:3]; // @[FlushableQueue.scala 33:24]
  wire [63:0] ram_instr__T_15_data; // @[FlushableQueue.scala 33:24]
  wire [1:0] ram_instr__T_15_addr; // @[FlushableQueue.scala 33:24]
  wire [63:0] ram_instr__T_5_data; // @[FlushableQueue.scala 33:24]
  wire [1:0] ram_instr__T_5_addr; // @[FlushableQueue.scala 33:24]
  wire  ram_instr__T_5_mask; // @[FlushableQueue.scala 33:24]
  wire  ram_instr__T_5_en; // @[FlushableQueue.scala 33:24]
  reg [38:0] ram_pc [0:3]; // @[FlushableQueue.scala 33:24]
  wire [38:0] ram_pc__T_15_data; // @[FlushableQueue.scala 33:24]
  wire [1:0] ram_pc__T_15_addr; // @[FlushableQueue.scala 33:24]
  wire [38:0] ram_pc__T_5_data; // @[FlushableQueue.scala 33:24]
  wire [1:0] ram_pc__T_5_addr; // @[FlushableQueue.scala 33:24]
  wire  ram_pc__T_5_mask; // @[FlushableQueue.scala 33:24]
  wire  ram_pc__T_5_en; // @[FlushableQueue.scala 33:24]
  reg [38:0] ram_pnpc [0:3]; // @[FlushableQueue.scala 33:24]
  wire [38:0] ram_pnpc__T_15_data; // @[FlushableQueue.scala 33:24]
  wire [1:0] ram_pnpc__T_15_addr; // @[FlushableQueue.scala 33:24]
  wire [38:0] ram_pnpc__T_5_data; // @[FlushableQueue.scala 33:24]
  wire [1:0] ram_pnpc__T_5_addr; // @[FlushableQueue.scala 33:24]
  wire  ram_pnpc__T_5_mask; // @[FlushableQueue.scala 33:24]
  wire  ram_pnpc__T_5_en; // @[FlushableQueue.scala 33:24]
  reg  ram_exceptionVec_12 [0:3]; // @[FlushableQueue.scala 33:24]
  wire  ram_exceptionVec_12__T_15_data; // @[FlushableQueue.scala 33:24]
  wire [1:0] ram_exceptionVec_12__T_15_addr; // @[FlushableQueue.scala 33:24]
  wire  ram_exceptionVec_12__T_5_data; // @[FlushableQueue.scala 33:24]
  wire [1:0] ram_exceptionVec_12__T_5_addr; // @[FlushableQueue.scala 33:24]
  wire  ram_exceptionVec_12__T_5_mask; // @[FlushableQueue.scala 33:24]
  wire  ram_exceptionVec_12__T_5_en; // @[FlushableQueue.scala 33:24]
  reg [3:0] ram_brIdx [0:3]; // @[FlushableQueue.scala 33:24]
  wire [3:0] ram_brIdx__T_15_data; // @[FlushableQueue.scala 33:24]
  wire [1:0] ram_brIdx__T_15_addr; // @[FlushableQueue.scala 33:24]
  wire [3:0] ram_brIdx__T_5_data; // @[FlushableQueue.scala 33:24]
  wire [1:0] ram_brIdx__T_5_addr; // @[FlushableQueue.scala 33:24]
  wire  ram_brIdx__T_5_mask; // @[FlushableQueue.scala 33:24]
  wire  ram_brIdx__T_5_en; // @[FlushableQueue.scala 33:24]
  reg [1:0] value; // @[Counter.scala 29:33]
  reg [1:0] value_1; // @[Counter.scala 29:33]
  reg  maybe_full; // @[FlushableQueue.scala 36:35]
  wire  _T = value == value_1; // @[FlushableQueue.scala 38:41]
  wire  _T_1 = ~maybe_full; // @[FlushableQueue.scala 39:36]
  wire  empty = _T & _T_1; // @[FlushableQueue.scala 39:33]
  wire  _T_2 = _T & maybe_full; // @[FlushableQueue.scala 40:32]
  wire  do_enq = io_enq_ready & io_enq_valid; // @[Decoupled.scala 40:37]
  wire  do_deq = io_deq_ready & io_deq_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _T_8 = value + 2'h1; // @[Counter.scala 39:22]
  wire [1:0] _T_11 = value_1 + 2'h1; // @[Counter.scala 39:22]
  wire  _T_12 = do_enq != do_deq; // @[FlushableQueue.scala 51:16]
  assign ram_instr__T_15_addr = value_1;
  assign ram_instr__T_15_data = ram_instr[ram_instr__T_15_addr]; // @[FlushableQueue.scala 33:24]
  assign ram_instr__T_5_data = io_enq_bits_instr;
  assign ram_instr__T_5_addr = value;
  assign ram_instr__T_5_mask = 1'h1;
  assign ram_instr__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_pc__T_15_addr = value_1;
  assign ram_pc__T_15_data = ram_pc[ram_pc__T_15_addr]; // @[FlushableQueue.scala 33:24]
  assign ram_pc__T_5_data = io_enq_bits_pc;
  assign ram_pc__T_5_addr = value;
  assign ram_pc__T_5_mask = 1'h1;
  assign ram_pc__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_pnpc__T_15_addr = value_1;
  assign ram_pnpc__T_15_data = ram_pnpc[ram_pnpc__T_15_addr]; // @[FlushableQueue.scala 33:24]
  assign ram_pnpc__T_5_data = io_enq_bits_pnpc;
  assign ram_pnpc__T_5_addr = value;
  assign ram_pnpc__T_5_mask = 1'h1;
  assign ram_pnpc__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_exceptionVec_12__T_15_addr = value_1;
  assign ram_exceptionVec_12__T_15_data = ram_exceptionVec_12[ram_exceptionVec_12__T_15_addr]; // @[FlushableQueue.scala 33:24]
  assign ram_exceptionVec_12__T_5_data = io_enq_bits_exceptionVec_12;
  assign ram_exceptionVec_12__T_5_addr = value;
  assign ram_exceptionVec_12__T_5_mask = 1'h1;
  assign ram_exceptionVec_12__T_5_en = io_enq_ready & io_enq_valid;
  assign ram_brIdx__T_15_addr = value_1;
  assign ram_brIdx__T_15_data = ram_brIdx[ram_brIdx__T_15_addr]; // @[FlushableQueue.scala 33:24]
  assign ram_brIdx__T_5_data = io_enq_bits_brIdx;
  assign ram_brIdx__T_5_addr = value;
  assign ram_brIdx__T_5_mask = 1'h1;
  assign ram_brIdx__T_5_en = io_enq_ready & io_enq_valid;
  assign io_enq_ready = ~_T_2; // @[FlushableQueue.scala 56:16]
  assign io_deq_valid = ~empty; // @[FlushableQueue.scala 55:16]
  assign io_deq_bits_instr = ram_instr__T_15_data; // @[FlushableQueue.scala 57:15]
  assign io_deq_bits_pc = ram_pc__T_15_data; // @[FlushableQueue.scala 57:15]
  assign io_deq_bits_pnpc = ram_pnpc__T_15_data; // @[FlushableQueue.scala 57:15]
  assign io_deq_bits_exceptionVec_12 = ram_exceptionVec_12__T_15_data; // @[FlushableQueue.scala 57:15]
  assign io_deq_bits_brIdx = ram_brIdx__T_15_data; // @[FlushableQueue.scala 57:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_instr[initvar] = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_pc[initvar] = _RAND_1[38:0];
  _RAND_2 = {2{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_pnpc[initvar] = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_exceptionVec_12[initvar] = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 4; initvar = initvar+1)
    ram_brIdx[initvar] = _RAND_4[3:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  value = _RAND_5[1:0];
  _RAND_6 = {1{`RANDOM}};
  value_1 = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  maybe_full = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(ram_instr__T_5_en & ram_instr__T_5_mask) begin
      ram_instr[ram_instr__T_5_addr] <= ram_instr__T_5_data; // @[FlushableQueue.scala 33:24]
    end
    if(ram_pc__T_5_en & ram_pc__T_5_mask) begin
      ram_pc[ram_pc__T_5_addr] <= ram_pc__T_5_data; // @[FlushableQueue.scala 33:24]
    end
    if(ram_pnpc__T_5_en & ram_pnpc__T_5_mask) begin
      ram_pnpc[ram_pnpc__T_5_addr] <= ram_pnpc__T_5_data; // @[FlushableQueue.scala 33:24]
    end
    if(ram_exceptionVec_12__T_5_en & ram_exceptionVec_12__T_5_mask) begin
      ram_exceptionVec_12[ram_exceptionVec_12__T_5_addr] <= ram_exceptionVec_12__T_5_data; // @[FlushableQueue.scala 33:24]
    end
    if(ram_brIdx__T_5_en & ram_brIdx__T_5_mask) begin
      ram_brIdx[ram_brIdx__T_5_addr] <= ram_brIdx__T_5_data; // @[FlushableQueue.scala 33:24]
    end
    if (reset) begin
      value <= 2'h0;
    end else if (io_flush) begin
      value <= 2'h0;
    end else if (do_enq) begin
      value <= _T_8;
    end
    if (reset) begin
      value_1 <= 2'h0;
    end else if (io_flush) begin
      value_1 <= 2'h0;
    end else if (do_deq) begin
      value_1 <= _T_11;
    end
    if (reset) begin
      maybe_full <= 1'h0;
    end else if (io_flush) begin
      maybe_full <= 1'h0;
    end else if (_T_12) begin
      maybe_full <= do_enq;
    end
  end
endmodule
module Frontend_inorder(
  input         clock,
  input         reset,
  input         io_out_0_ready,
  output        io_out_0_valid,
  output [63:0] io_out_0_bits_cf_instr,
  output [38:0] io_out_0_bits_cf_pc,
  output [38:0] io_out_0_bits_cf_pnpc,
  output        io_out_0_bits_cf_exceptionVec_1,
  output        io_out_0_bits_cf_exceptionVec_2,
  output        io_out_0_bits_cf_exceptionVec_12,
  output        io_out_0_bits_cf_intrVec_0,
  output        io_out_0_bits_cf_intrVec_1,
  output        io_out_0_bits_cf_intrVec_2,
  output        io_out_0_bits_cf_intrVec_3,
  output        io_out_0_bits_cf_intrVec_4,
  output        io_out_0_bits_cf_intrVec_5,
  output        io_out_0_bits_cf_intrVec_6,
  output        io_out_0_bits_cf_intrVec_7,
  output        io_out_0_bits_cf_intrVec_8,
  output        io_out_0_bits_cf_intrVec_9,
  output        io_out_0_bits_cf_intrVec_10,
  output        io_out_0_bits_cf_intrVec_11,
  output [3:0]  io_out_0_bits_cf_brIdx,
  output        io_out_0_bits_cf_crossPageIPFFix,
  output        io_out_0_bits_ctrl_src1Type,
  output        io_out_0_bits_ctrl_src2Type,
  output [2:0]  io_out_0_bits_ctrl_fuType,
  output [6:0]  io_out_0_bits_ctrl_fuOpType,
  output [4:0]  io_out_0_bits_ctrl_rfSrc1,
  output [4:0]  io_out_0_bits_ctrl_rfSrc2,
  output        io_out_0_bits_ctrl_rfWen,
  output [4:0]  io_out_0_bits_ctrl_rfDest,
  output [63:0] io_out_0_bits_data_imm,
  output        io_out_1_bits_cf_intrVec_0,
  output        io_out_1_bits_cf_intrVec_1,
  output        io_out_1_bits_cf_intrVec_2,
  output        io_out_1_bits_cf_intrVec_3,
  output        io_out_1_bits_cf_intrVec_4,
  output        io_out_1_bits_cf_intrVec_5,
  output        io_out_1_bits_cf_intrVec_6,
  output        io_out_1_bits_cf_intrVec_7,
  output        io_out_1_bits_cf_intrVec_8,
  output        io_out_1_bits_cf_intrVec_9,
  output        io_out_1_bits_cf_intrVec_10,
  output        io_out_1_bits_cf_intrVec_11,
  input         io_imem_req_ready,
  output        io_imem_req_valid,
  output [38:0] io_imem_req_bits_addr,
  output [86:0] io_imem_req_bits_user,
  output        io_imem_resp_ready,
  input         io_imem_resp_valid,
  input  [63:0] io_imem_resp_bits_rdata,
  input  [86:0] io_imem_resp_bits_user,
  output [3:0]  io_flushVec,
  input         io_ipf,
  input  [38:0] io_redirect_target,
  input         io_redirect_valid,
  input         flushICache,
  input         _T_243_valid,
  input  [38:0] _T_243_pc,
  input         _T_243_isMissPredict,
  input  [38:0] _T_243_actualTarget,
  input         _T_243_actualTaken,
  input  [6:0]  _T_243_fuOpType,
  input  [1:0]  _T_243_btbType,
  input         _T_243_isRVC,
  input         vmEnable,
  input  [11:0] intrVec,
  input         flushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  ifu_clock; // @[Frontend.scala 106:20]
  wire  ifu_reset; // @[Frontend.scala 106:20]
  wire  ifu_io_imem_req_ready; // @[Frontend.scala 106:20]
  wire  ifu_io_imem_req_valid; // @[Frontend.scala 106:20]
  wire [38:0] ifu_io_imem_req_bits_addr; // @[Frontend.scala 106:20]
  wire [81:0] ifu_io_imem_req_bits_user; // @[Frontend.scala 106:20]
  wire  ifu_io_imem_resp_ready; // @[Frontend.scala 106:20]
  wire  ifu_io_imem_resp_valid; // @[Frontend.scala 106:20]
  wire [63:0] ifu_io_imem_resp_bits_rdata; // @[Frontend.scala 106:20]
  wire [81:0] ifu_io_imem_resp_bits_user; // @[Frontend.scala 106:20]
  wire  ifu_io_out_ready; // @[Frontend.scala 106:20]
  wire  ifu_io_out_valid; // @[Frontend.scala 106:20]
  wire [63:0] ifu_io_out_bits_instr; // @[Frontend.scala 106:20]
  wire [38:0] ifu_io_out_bits_pc; // @[Frontend.scala 106:20]
  wire [38:0] ifu_io_out_bits_pnpc; // @[Frontend.scala 106:20]
  wire  ifu_io_out_bits_exceptionVec_12; // @[Frontend.scala 106:20]
  wire [3:0] ifu_io_out_bits_brIdx; // @[Frontend.scala 106:20]
  wire [38:0] ifu_io_redirect_target; // @[Frontend.scala 106:20]
  wire  ifu_io_redirect_valid; // @[Frontend.scala 106:20]
  wire [3:0] ifu_io_flushVec; // @[Frontend.scala 106:20]
  wire  ifu_io_ipf; // @[Frontend.scala 106:20]
  wire  ifu_flushICache; // @[Frontend.scala 106:20]
  wire  ifu__T_243_valid; // @[Frontend.scala 106:20]
  wire [38:0] ifu__T_243_pc; // @[Frontend.scala 106:20]
  wire  ifu__T_243_isMissPredict; // @[Frontend.scala 106:20]
  wire [38:0] ifu__T_243_actualTarget; // @[Frontend.scala 106:20]
  wire  ifu__T_243_actualTaken; // @[Frontend.scala 106:20]
  wire [6:0] ifu__T_243_fuOpType; // @[Frontend.scala 106:20]
  wire [1:0] ifu__T_243_btbType; // @[Frontend.scala 106:20]
  wire  ifu__T_243_isRVC; // @[Frontend.scala 106:20]
  wire  ifu_flushTLB; // @[Frontend.scala 106:20]
  wire  ibf_clock; // @[Frontend.scala 107:19]
  wire  ibf_reset; // @[Frontend.scala 107:19]
  wire  ibf_io_in_ready; // @[Frontend.scala 107:19]
  wire  ibf_io_in_valid; // @[Frontend.scala 107:19]
  wire [63:0] ibf_io_in_bits_instr; // @[Frontend.scala 107:19]
  wire [38:0] ibf_io_in_bits_pc; // @[Frontend.scala 107:19]
  wire [38:0] ibf_io_in_bits_pnpc; // @[Frontend.scala 107:19]
  wire  ibf_io_in_bits_exceptionVec_12; // @[Frontend.scala 107:19]
  wire [3:0] ibf_io_in_bits_brIdx; // @[Frontend.scala 107:19]
  wire  ibf_io_out_ready; // @[Frontend.scala 107:19]
  wire  ibf_io_out_valid; // @[Frontend.scala 107:19]
  wire [63:0] ibf_io_out_bits_instr; // @[Frontend.scala 107:19]
  wire [38:0] ibf_io_out_bits_pc; // @[Frontend.scala 107:19]
  wire [38:0] ibf_io_out_bits_pnpc; // @[Frontend.scala 107:19]
  wire  ibf_io_out_bits_exceptionVec_12; // @[Frontend.scala 107:19]
  wire [3:0] ibf_io_out_bits_brIdx; // @[Frontend.scala 107:19]
  wire  ibf_io_out_bits_crossPageIPFFix; // @[Frontend.scala 107:19]
  wire  ibf_io_flush; // @[Frontend.scala 107:19]
  wire  idu_io_in_0_ready; // @[Frontend.scala 108:20]
  wire  idu_io_in_0_valid; // @[Frontend.scala 108:20]
  wire [63:0] idu_io_in_0_bits_instr; // @[Frontend.scala 108:20]
  wire [38:0] idu_io_in_0_bits_pc; // @[Frontend.scala 108:20]
  wire [38:0] idu_io_in_0_bits_pnpc; // @[Frontend.scala 108:20]
  wire  idu_io_in_0_bits_exceptionVec_12; // @[Frontend.scala 108:20]
  wire [3:0] idu_io_in_0_bits_brIdx; // @[Frontend.scala 108:20]
  wire  idu_io_in_0_bits_crossPageIPFFix; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_ready; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_valid; // @[Frontend.scala 108:20]
  wire [63:0] idu_io_out_0_bits_cf_instr; // @[Frontend.scala 108:20]
  wire [38:0] idu_io_out_0_bits_cf_pc; // @[Frontend.scala 108:20]
  wire [38:0] idu_io_out_0_bits_cf_pnpc; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_1; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_2; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_exceptionVec_12; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_0; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_1; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_2; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_3; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_4; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_5; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_6; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_7; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_8; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_9; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_10; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_intrVec_11; // @[Frontend.scala 108:20]
  wire [3:0] idu_io_out_0_bits_cf_brIdx; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_cf_crossPageIPFFix; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_ctrl_src1Type; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_ctrl_src2Type; // @[Frontend.scala 108:20]
  wire [2:0] idu_io_out_0_bits_ctrl_fuType; // @[Frontend.scala 108:20]
  wire [6:0] idu_io_out_0_bits_ctrl_fuOpType; // @[Frontend.scala 108:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfSrc1; // @[Frontend.scala 108:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfSrc2; // @[Frontend.scala 108:20]
  wire  idu_io_out_0_bits_ctrl_rfWen; // @[Frontend.scala 108:20]
  wire [4:0] idu_io_out_0_bits_ctrl_rfDest; // @[Frontend.scala 108:20]
  wire [63:0] idu_io_out_0_bits_data_imm; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_0; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_1; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_2; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_3; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_4; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_5; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_6; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_7; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_8; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_9; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_10; // @[Frontend.scala 108:20]
  wire  idu_io_out_1_bits_cf_intrVec_11; // @[Frontend.scala 108:20]
  wire  idu_vmEnable; // @[Frontend.scala 108:20]
  wire [11:0] idu_intrVec; // @[Frontend.scala 108:20]
  wire  FlushableQueue_clock; // @[FlushableQueue.scala 104:21]
  wire  FlushableQueue_reset; // @[FlushableQueue.scala 104:21]
  wire  FlushableQueue_io_enq_ready; // @[FlushableQueue.scala 104:21]
  wire  FlushableQueue_io_enq_valid; // @[FlushableQueue.scala 104:21]
  wire [63:0] FlushableQueue_io_enq_bits_instr; // @[FlushableQueue.scala 104:21]
  wire [38:0] FlushableQueue_io_enq_bits_pc; // @[FlushableQueue.scala 104:21]
  wire [38:0] FlushableQueue_io_enq_bits_pnpc; // @[FlushableQueue.scala 104:21]
  wire  FlushableQueue_io_enq_bits_exceptionVec_12; // @[FlushableQueue.scala 104:21]
  wire [3:0] FlushableQueue_io_enq_bits_brIdx; // @[FlushableQueue.scala 104:21]
  wire  FlushableQueue_io_deq_ready; // @[FlushableQueue.scala 104:21]
  wire  FlushableQueue_io_deq_valid; // @[FlushableQueue.scala 104:21]
  wire [63:0] FlushableQueue_io_deq_bits_instr; // @[FlushableQueue.scala 104:21]
  wire [38:0] FlushableQueue_io_deq_bits_pc; // @[FlushableQueue.scala 104:21]
  wire [38:0] FlushableQueue_io_deq_bits_pnpc; // @[FlushableQueue.scala 104:21]
  wire  FlushableQueue_io_deq_bits_exceptionVec_12; // @[FlushableQueue.scala 104:21]
  wire [3:0] FlushableQueue_io_deq_bits_brIdx; // @[FlushableQueue.scala 104:21]
  wire  FlushableQueue_io_flush; // @[FlushableQueue.scala 104:21]
  wire  _T_1 = idu_io_out_0_ready & idu_io_out_0_valid; // @[Decoupled.scala 40:37]
  reg  _T_3; // @[Pipeline.scala 24:24]
  wire  _GEN_0 = _T_1 ? 1'h0 : _T_3; // @[Pipeline.scala 25:25]
  wire  _T_4 = ibf_io_out_valid & idu_io_in_0_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_1 = _T_4 | _GEN_0; // @[Pipeline.scala 26:38]
  reg [63:0] _T_6_instr; // @[Reg.scala 15:16]
  reg [38:0] _T_6_pc; // @[Reg.scala 15:16]
  reg [38:0] _T_6_pnpc; // @[Reg.scala 15:16]
  reg  _T_6_exceptionVec_12; // @[Reg.scala 15:16]
  reg [3:0] _T_6_brIdx; // @[Reg.scala 15:16]
  reg  _T_6_crossPageIPFFix; // @[Reg.scala 15:16]
  IFU_inorder ifu ( // @[Frontend.scala 106:20]
    .clock(ifu_clock),
    .reset(ifu_reset),
    .io_imem_req_ready(ifu_io_imem_req_ready),
    .io_imem_req_valid(ifu_io_imem_req_valid),
    .io_imem_req_bits_addr(ifu_io_imem_req_bits_addr),
    .io_imem_req_bits_user(ifu_io_imem_req_bits_user),
    .io_imem_resp_ready(ifu_io_imem_resp_ready),
    .io_imem_resp_valid(ifu_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(ifu_io_imem_resp_bits_rdata),
    .io_imem_resp_bits_user(ifu_io_imem_resp_bits_user),
    .io_out_ready(ifu_io_out_ready),
    .io_out_valid(ifu_io_out_valid),
    .io_out_bits_instr(ifu_io_out_bits_instr),
    .io_out_bits_pc(ifu_io_out_bits_pc),
    .io_out_bits_pnpc(ifu_io_out_bits_pnpc),
    .io_out_bits_exceptionVec_12(ifu_io_out_bits_exceptionVec_12),
    .io_out_bits_brIdx(ifu_io_out_bits_brIdx),
    .io_redirect_target(ifu_io_redirect_target),
    .io_redirect_valid(ifu_io_redirect_valid),
    .io_flushVec(ifu_io_flushVec),
    .io_ipf(ifu_io_ipf),
    .flushICache(ifu_flushICache),
    ._T_243_valid(ifu__T_243_valid),
    ._T_243_pc(ifu__T_243_pc),
    ._T_243_isMissPredict(ifu__T_243_isMissPredict),
    ._T_243_actualTarget(ifu__T_243_actualTarget),
    ._T_243_actualTaken(ifu__T_243_actualTaken),
    ._T_243_fuOpType(ifu__T_243_fuOpType),
    ._T_243_btbType(ifu__T_243_btbType),
    ._T_243_isRVC(ifu__T_243_isRVC),
    .flushTLB(ifu_flushTLB)
  );
  NaiveRVCAlignBuffer ibf ( // @[Frontend.scala 107:19]
    .clock(ibf_clock),
    .reset(ibf_reset),
    .io_in_ready(ibf_io_in_ready),
    .io_in_valid(ibf_io_in_valid),
    .io_in_bits_instr(ibf_io_in_bits_instr),
    .io_in_bits_pc(ibf_io_in_bits_pc),
    .io_in_bits_pnpc(ibf_io_in_bits_pnpc),
    .io_in_bits_exceptionVec_12(ibf_io_in_bits_exceptionVec_12),
    .io_in_bits_brIdx(ibf_io_in_bits_brIdx),
    .io_out_ready(ibf_io_out_ready),
    .io_out_valid(ibf_io_out_valid),
    .io_out_bits_instr(ibf_io_out_bits_instr),
    .io_out_bits_pc(ibf_io_out_bits_pc),
    .io_out_bits_pnpc(ibf_io_out_bits_pnpc),
    .io_out_bits_exceptionVec_12(ibf_io_out_bits_exceptionVec_12),
    .io_out_bits_brIdx(ibf_io_out_bits_brIdx),
    .io_out_bits_crossPageIPFFix(ibf_io_out_bits_crossPageIPFFix),
    .io_flush(ibf_io_flush)
  );
  IDU idu ( // @[Frontend.scala 108:20]
    .io_in_0_ready(idu_io_in_0_ready),
    .io_in_0_valid(idu_io_in_0_valid),
    .io_in_0_bits_instr(idu_io_in_0_bits_instr),
    .io_in_0_bits_pc(idu_io_in_0_bits_pc),
    .io_in_0_bits_pnpc(idu_io_in_0_bits_pnpc),
    .io_in_0_bits_exceptionVec_12(idu_io_in_0_bits_exceptionVec_12),
    .io_in_0_bits_brIdx(idu_io_in_0_bits_brIdx),
    .io_in_0_bits_crossPageIPFFix(idu_io_in_0_bits_crossPageIPFFix),
    .io_out_0_ready(idu_io_out_0_ready),
    .io_out_0_valid(idu_io_out_0_valid),
    .io_out_0_bits_cf_instr(idu_io_out_0_bits_cf_instr),
    .io_out_0_bits_cf_pc(idu_io_out_0_bits_cf_pc),
    .io_out_0_bits_cf_pnpc(idu_io_out_0_bits_cf_pnpc),
    .io_out_0_bits_cf_exceptionVec_1(idu_io_out_0_bits_cf_exceptionVec_1),
    .io_out_0_bits_cf_exceptionVec_2(idu_io_out_0_bits_cf_exceptionVec_2),
    .io_out_0_bits_cf_exceptionVec_12(idu_io_out_0_bits_cf_exceptionVec_12),
    .io_out_0_bits_cf_intrVec_0(idu_io_out_0_bits_cf_intrVec_0),
    .io_out_0_bits_cf_intrVec_1(idu_io_out_0_bits_cf_intrVec_1),
    .io_out_0_bits_cf_intrVec_2(idu_io_out_0_bits_cf_intrVec_2),
    .io_out_0_bits_cf_intrVec_3(idu_io_out_0_bits_cf_intrVec_3),
    .io_out_0_bits_cf_intrVec_4(idu_io_out_0_bits_cf_intrVec_4),
    .io_out_0_bits_cf_intrVec_5(idu_io_out_0_bits_cf_intrVec_5),
    .io_out_0_bits_cf_intrVec_6(idu_io_out_0_bits_cf_intrVec_6),
    .io_out_0_bits_cf_intrVec_7(idu_io_out_0_bits_cf_intrVec_7),
    .io_out_0_bits_cf_intrVec_8(idu_io_out_0_bits_cf_intrVec_8),
    .io_out_0_bits_cf_intrVec_9(idu_io_out_0_bits_cf_intrVec_9),
    .io_out_0_bits_cf_intrVec_10(idu_io_out_0_bits_cf_intrVec_10),
    .io_out_0_bits_cf_intrVec_11(idu_io_out_0_bits_cf_intrVec_11),
    .io_out_0_bits_cf_brIdx(idu_io_out_0_bits_cf_brIdx),
    .io_out_0_bits_cf_crossPageIPFFix(idu_io_out_0_bits_cf_crossPageIPFFix),
    .io_out_0_bits_ctrl_src1Type(idu_io_out_0_bits_ctrl_src1Type),
    .io_out_0_bits_ctrl_src2Type(idu_io_out_0_bits_ctrl_src2Type),
    .io_out_0_bits_ctrl_fuType(idu_io_out_0_bits_ctrl_fuType),
    .io_out_0_bits_ctrl_fuOpType(idu_io_out_0_bits_ctrl_fuOpType),
    .io_out_0_bits_ctrl_rfSrc1(idu_io_out_0_bits_ctrl_rfSrc1),
    .io_out_0_bits_ctrl_rfSrc2(idu_io_out_0_bits_ctrl_rfSrc2),
    .io_out_0_bits_ctrl_rfWen(idu_io_out_0_bits_ctrl_rfWen),
    .io_out_0_bits_ctrl_rfDest(idu_io_out_0_bits_ctrl_rfDest),
    .io_out_0_bits_data_imm(idu_io_out_0_bits_data_imm),
    .io_out_1_bits_cf_intrVec_0(idu_io_out_1_bits_cf_intrVec_0),
    .io_out_1_bits_cf_intrVec_1(idu_io_out_1_bits_cf_intrVec_1),
    .io_out_1_bits_cf_intrVec_2(idu_io_out_1_bits_cf_intrVec_2),
    .io_out_1_bits_cf_intrVec_3(idu_io_out_1_bits_cf_intrVec_3),
    .io_out_1_bits_cf_intrVec_4(idu_io_out_1_bits_cf_intrVec_4),
    .io_out_1_bits_cf_intrVec_5(idu_io_out_1_bits_cf_intrVec_5),
    .io_out_1_bits_cf_intrVec_6(idu_io_out_1_bits_cf_intrVec_6),
    .io_out_1_bits_cf_intrVec_7(idu_io_out_1_bits_cf_intrVec_7),
    .io_out_1_bits_cf_intrVec_8(idu_io_out_1_bits_cf_intrVec_8),
    .io_out_1_bits_cf_intrVec_9(idu_io_out_1_bits_cf_intrVec_9),
    .io_out_1_bits_cf_intrVec_10(idu_io_out_1_bits_cf_intrVec_10),
    .io_out_1_bits_cf_intrVec_11(idu_io_out_1_bits_cf_intrVec_11),
    .vmEnable(idu_vmEnable),
    .intrVec(idu_intrVec)
  );
  FlushableQueue FlushableQueue ( // @[FlushableQueue.scala 104:21]
    .clock(FlushableQueue_clock),
    .reset(FlushableQueue_reset),
    .io_enq_ready(FlushableQueue_io_enq_ready),
    .io_enq_valid(FlushableQueue_io_enq_valid),
    .io_enq_bits_instr(FlushableQueue_io_enq_bits_instr),
    .io_enq_bits_pc(FlushableQueue_io_enq_bits_pc),
    .io_enq_bits_pnpc(FlushableQueue_io_enq_bits_pnpc),
    .io_enq_bits_exceptionVec_12(FlushableQueue_io_enq_bits_exceptionVec_12),
    .io_enq_bits_brIdx(FlushableQueue_io_enq_bits_brIdx),
    .io_deq_ready(FlushableQueue_io_deq_ready),
    .io_deq_valid(FlushableQueue_io_deq_valid),
    .io_deq_bits_instr(FlushableQueue_io_deq_bits_instr),
    .io_deq_bits_pc(FlushableQueue_io_deq_bits_pc),
    .io_deq_bits_pnpc(FlushableQueue_io_deq_bits_pnpc),
    .io_deq_bits_exceptionVec_12(FlushableQueue_io_deq_bits_exceptionVec_12),
    .io_deq_bits_brIdx(FlushableQueue_io_deq_bits_brIdx),
    .io_flush(FlushableQueue_io_flush)
  );
  assign io_out_0_valid = idu_io_out_0_valid; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_instr = idu_io_out_0_bits_cf_instr; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_pc = idu_io_out_0_bits_cf_pc; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_pnpc = idu_io_out_0_bits_cf_pnpc; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_exceptionVec_1 = idu_io_out_0_bits_cf_exceptionVec_1; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_exceptionVec_2 = idu_io_out_0_bits_cf_exceptionVec_2; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_exceptionVec_12 = idu_io_out_0_bits_cf_exceptionVec_12; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_0 = idu_io_out_0_bits_cf_intrVec_0; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_1 = idu_io_out_0_bits_cf_intrVec_1; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_2 = idu_io_out_0_bits_cf_intrVec_2; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_3 = idu_io_out_0_bits_cf_intrVec_3; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_4 = idu_io_out_0_bits_cf_intrVec_4; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_5 = idu_io_out_0_bits_cf_intrVec_5; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_6 = idu_io_out_0_bits_cf_intrVec_6; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_7 = idu_io_out_0_bits_cf_intrVec_7; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_8 = idu_io_out_0_bits_cf_intrVec_8; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_9 = idu_io_out_0_bits_cf_intrVec_9; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_10 = idu_io_out_0_bits_cf_intrVec_10; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_intrVec_11 = idu_io_out_0_bits_cf_intrVec_11; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_brIdx = idu_io_out_0_bits_cf_brIdx; // @[Frontend.scala 120:10]
  assign io_out_0_bits_cf_crossPageIPFFix = idu_io_out_0_bits_cf_crossPageIPFFix; // @[Frontend.scala 120:10]
  assign io_out_0_bits_ctrl_src1Type = idu_io_out_0_bits_ctrl_src1Type; // @[Frontend.scala 120:10]
  assign io_out_0_bits_ctrl_src2Type = idu_io_out_0_bits_ctrl_src2Type; // @[Frontend.scala 120:10]
  assign io_out_0_bits_ctrl_fuType = idu_io_out_0_bits_ctrl_fuType; // @[Frontend.scala 120:10]
  assign io_out_0_bits_ctrl_fuOpType = idu_io_out_0_bits_ctrl_fuOpType; // @[Frontend.scala 120:10]
  assign io_out_0_bits_ctrl_rfSrc1 = idu_io_out_0_bits_ctrl_rfSrc1; // @[Frontend.scala 120:10]
  assign io_out_0_bits_ctrl_rfSrc2 = idu_io_out_0_bits_ctrl_rfSrc2; // @[Frontend.scala 120:10]
  assign io_out_0_bits_ctrl_rfWen = idu_io_out_0_bits_ctrl_rfWen; // @[Frontend.scala 120:10]
  assign io_out_0_bits_ctrl_rfDest = idu_io_out_0_bits_ctrl_rfDest; // @[Frontend.scala 120:10]
  assign io_out_0_bits_data_imm = idu_io_out_0_bits_data_imm; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_0 = idu_io_out_1_bits_cf_intrVec_0; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_1 = idu_io_out_1_bits_cf_intrVec_1; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_2 = idu_io_out_1_bits_cf_intrVec_2; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_3 = idu_io_out_1_bits_cf_intrVec_3; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_4 = idu_io_out_1_bits_cf_intrVec_4; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_5 = idu_io_out_1_bits_cf_intrVec_5; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_6 = idu_io_out_1_bits_cf_intrVec_6; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_7 = idu_io_out_1_bits_cf_intrVec_7; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_8 = idu_io_out_1_bits_cf_intrVec_8; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_9 = idu_io_out_1_bits_cf_intrVec_9; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_10 = idu_io_out_1_bits_cf_intrVec_10; // @[Frontend.scala 120:10]
  assign io_out_1_bits_cf_intrVec_11 = idu_io_out_1_bits_cf_intrVec_11; // @[Frontend.scala 120:10]
  assign io_imem_req_valid = ifu_io_imem_req_valid; // @[Frontend.scala 125:11]
  assign io_imem_req_bits_addr = ifu_io_imem_req_bits_addr; // @[Frontend.scala 125:11]
  assign io_imem_req_bits_user = {{5'd0}, ifu_io_imem_req_bits_user}; // @[Frontend.scala 125:11]
  assign io_imem_resp_ready = ifu_io_imem_resp_ready; // @[Frontend.scala 125:11]
  assign io_flushVec = ifu_io_flushVec; // @[Frontend.scala 122:15]
  assign ifu_clock = clock;
  assign ifu_reset = reset;
  assign ifu_io_imem_req_ready = io_imem_req_ready; // @[Frontend.scala 125:11]
  assign ifu_io_imem_resp_valid = io_imem_resp_valid; // @[Frontend.scala 125:11]
  assign ifu_io_imem_resp_bits_rdata = io_imem_resp_bits_rdata; // @[Frontend.scala 125:11]
  assign ifu_io_imem_resp_bits_user = io_imem_resp_bits_user[81:0]; // @[Frontend.scala 125:11]
  assign ifu_io_out_ready = FlushableQueue_io_enq_ready; // @[FlushableQueue.scala 108:17]
  assign ifu_io_redirect_target = io_redirect_target; // @[Frontend.scala 121:15]
  assign ifu_io_redirect_valid = io_redirect_valid; // @[Frontend.scala 121:15]
  assign ifu_io_ipf = io_ipf; // @[Frontend.scala 124:10]
  assign ifu_flushICache = flushICache;
  assign ifu__T_243_valid = _T_243_valid;
  assign ifu__T_243_pc = _T_243_pc;
  assign ifu__T_243_isMissPredict = _T_243_isMissPredict;
  assign ifu__T_243_actualTarget = _T_243_actualTarget;
  assign ifu__T_243_actualTaken = _T_243_actualTaken;
  assign ifu__T_243_fuOpType = _T_243_fuOpType;
  assign ifu__T_243_btbType = _T_243_btbType;
  assign ifu__T_243_isRVC = _T_243_isRVC;
  assign ifu_flushTLB = flushTLB;
  assign ibf_clock = clock;
  assign ibf_reset = reset;
  assign ibf_io_in_valid = FlushableQueue_io_deq_valid; // @[Frontend.scala 112:11]
  assign ibf_io_in_bits_instr = FlushableQueue_io_deq_bits_instr; // @[Frontend.scala 112:11]
  assign ibf_io_in_bits_pc = FlushableQueue_io_deq_bits_pc; // @[Frontend.scala 112:11]
  assign ibf_io_in_bits_pnpc = FlushableQueue_io_deq_bits_pnpc; // @[Frontend.scala 112:11]
  assign ibf_io_in_bits_exceptionVec_12 = FlushableQueue_io_deq_bits_exceptionVec_12; // @[Frontend.scala 112:11]
  assign ibf_io_in_bits_brIdx = FlushableQueue_io_deq_bits_brIdx; // @[Frontend.scala 112:11]
  assign ibf_io_out_ready = idu_io_in_0_ready; // @[Pipeline.scala 29:16]
  assign ibf_io_flush = ifu_io_flushVec[1]; // @[Frontend.scala 119:16]
  assign idu_io_in_0_valid = _T_3; // @[Pipeline.scala 31:17]
  assign idu_io_in_0_bits_instr = _T_6_instr; // @[Pipeline.scala 30:16]
  assign idu_io_in_0_bits_pc = _T_6_pc; // @[Pipeline.scala 30:16]
  assign idu_io_in_0_bits_pnpc = _T_6_pnpc; // @[Pipeline.scala 30:16]
  assign idu_io_in_0_bits_exceptionVec_12 = _T_6_exceptionVec_12; // @[Pipeline.scala 30:16]
  assign idu_io_in_0_bits_brIdx = _T_6_brIdx; // @[Pipeline.scala 30:16]
  assign idu_io_in_0_bits_crossPageIPFFix = _T_6_crossPageIPFFix; // @[Pipeline.scala 30:16]
  assign idu_io_out_0_ready = io_out_0_ready; // @[Frontend.scala 120:10]
  assign idu_vmEnable = vmEnable;
  assign idu_intrVec = intrVec;
  assign FlushableQueue_clock = clock;
  assign FlushableQueue_reset = reset;
  assign FlushableQueue_io_enq_valid = ifu_io_out_valid; // @[FlushableQueue.scala 105:22]
  assign FlushableQueue_io_enq_bits_instr = ifu_io_out_bits_instr; // @[FlushableQueue.scala 106:21]
  assign FlushableQueue_io_enq_bits_pc = ifu_io_out_bits_pc; // @[FlushableQueue.scala 106:21]
  assign FlushableQueue_io_enq_bits_pnpc = ifu_io_out_bits_pnpc; // @[FlushableQueue.scala 106:21]
  assign FlushableQueue_io_enq_bits_exceptionVec_12 = ifu_io_out_bits_exceptionVec_12; // @[FlushableQueue.scala 106:21]
  assign FlushableQueue_io_enq_bits_brIdx = ifu_io_out_bits_brIdx; // @[FlushableQueue.scala 106:21]
  assign FlushableQueue_io_deq_ready = ibf_io_in_ready; // @[Frontend.scala 112:11]
  assign FlushableQueue_io_flush = ifu_io_flushVec[0]; // @[FlushableQueue.scala 107:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_3 = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  _T_6_instr = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  _T_6_pc = _RAND_2[38:0];
  _RAND_3 = {2{`RANDOM}};
  _T_6_pnpc = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  _T_6_exceptionVec_12 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_6_brIdx = _RAND_5[3:0];
  _RAND_6 = {1{`RANDOM}};
  _T_6_crossPageIPFFix = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_3 <= 1'h0;
    end else if (ifu_io_flushVec[1]) begin
      _T_3 <= 1'h0;
    end else begin
      _T_3 <= _GEN_1;
    end
    if (_T_4) begin
      _T_6_instr <= ibf_io_out_bits_instr;
    end
    if (_T_4) begin
      _T_6_pc <= ibf_io_out_bits_pc;
    end
    if (_T_4) begin
      _T_6_pnpc <= ibf_io_out_bits_pnpc;
    end
    if (_T_4) begin
      _T_6_exceptionVec_12 <= ibf_io_out_bits_exceptionVec_12;
    end
    if (_T_4) begin
      _T_6_brIdx <= ibf_io_out_bits_brIdx;
    end
    if (_T_4) begin
      _T_6_crossPageIPFFix <= ibf_io_out_bits_crossPageIPFFix;
    end
  end
endmodule
module ISU(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [63:0] io_in_0_bits_cf_instr,
  input  [38:0] io_in_0_bits_cf_pc,
  input  [38:0] io_in_0_bits_cf_pnpc,
  input         io_in_0_bits_cf_exceptionVec_1,
  input         io_in_0_bits_cf_exceptionVec_2,
  input         io_in_0_bits_cf_exceptionVec_12,
  input         io_in_0_bits_cf_intrVec_0,
  input         io_in_0_bits_cf_intrVec_1,
  input         io_in_0_bits_cf_intrVec_2,
  input         io_in_0_bits_cf_intrVec_3,
  input         io_in_0_bits_cf_intrVec_4,
  input         io_in_0_bits_cf_intrVec_5,
  input         io_in_0_bits_cf_intrVec_6,
  input         io_in_0_bits_cf_intrVec_7,
  input         io_in_0_bits_cf_intrVec_8,
  input         io_in_0_bits_cf_intrVec_9,
  input         io_in_0_bits_cf_intrVec_10,
  input         io_in_0_bits_cf_intrVec_11,
  input  [3:0]  io_in_0_bits_cf_brIdx,
  input         io_in_0_bits_cf_crossPageIPFFix,
  input         io_in_0_bits_ctrl_src1Type,
  input         io_in_0_bits_ctrl_src2Type,
  input  [2:0]  io_in_0_bits_ctrl_fuType,
  input  [6:0]  io_in_0_bits_ctrl_fuOpType,
  input  [4:0]  io_in_0_bits_ctrl_rfSrc1,
  input  [4:0]  io_in_0_bits_ctrl_rfSrc2,
  input         io_in_0_bits_ctrl_rfWen,
  input  [4:0]  io_in_0_bits_ctrl_rfDest,
  input  [63:0] io_in_0_bits_data_imm,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_cf_instr,
  output [38:0] io_out_bits_cf_pc,
  output [38:0] io_out_bits_cf_pnpc,
  output        io_out_bits_cf_exceptionVec_1,
  output        io_out_bits_cf_exceptionVec_2,
  output        io_out_bits_cf_exceptionVec_12,
  output        io_out_bits_cf_intrVec_0,
  output        io_out_bits_cf_intrVec_1,
  output        io_out_bits_cf_intrVec_2,
  output        io_out_bits_cf_intrVec_3,
  output        io_out_bits_cf_intrVec_4,
  output        io_out_bits_cf_intrVec_5,
  output        io_out_bits_cf_intrVec_6,
  output        io_out_bits_cf_intrVec_7,
  output        io_out_bits_cf_intrVec_8,
  output        io_out_bits_cf_intrVec_9,
  output        io_out_bits_cf_intrVec_10,
  output        io_out_bits_cf_intrVec_11,
  output [3:0]  io_out_bits_cf_brIdx,
  output        io_out_bits_cf_crossPageIPFFix,
  output [2:0]  io_out_bits_ctrl_fuType,
  output [6:0]  io_out_bits_ctrl_fuOpType,
  output        io_out_bits_ctrl_rfWen,
  output [4:0]  io_out_bits_ctrl_rfDest,
  output [63:0] io_out_bits_data_src1,
  output [63:0] io_out_bits_data_src2,
  output [63:0] io_out_bits_data_imm,
  input         io_wb_rfWen,
  input  [4:0]  io_wb_rfDest,
  input  [63:0] io_wb_rfData,
  input         io_forward_valid,
  input         io_forward_wb_rfWen,
  input  [4:0]  io_forward_wb_rfDest,
  input  [63:0] io_forward_wb_rfData,
  input  [2:0]  io_forward_fuType,
  input         io_flush
);
`ifdef RANDOMIZE_MEM_INIT
  reg [63:0] _RAND_0;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] _T_31 [0:31]; // @[RF.scala 30:15]
  wire [63:0] _T_31__T_45_data; // @[RF.scala 30:15]
  wire [4:0] _T_31__T_45_addr; // @[RF.scala 30:15]
  wire [63:0] _T_31__T_64_data; // @[RF.scala 30:15]
  wire [4:0] _T_31__T_64_addr; // @[RF.scala 30:15]
  wire [63:0] _T_31__T_74_data; // @[RF.scala 30:15]
  wire [4:0] _T_31__T_74_addr; // @[RF.scala 30:15]
  wire  _T_31__T_74_mask; // @[RF.scala 30:15]
  wire  _T_31__T_74_en; // @[RF.scala 30:15]
  wire  forwardRfWen = io_forward_wb_rfWen & io_forward_valid; // @[ISU.scala 42:42]
  wire  _T = io_forward_fuType != 3'h0; // @[ISU.scala 43:41]
  wire  _T_1 = io_forward_fuType != 3'h1; // @[ISU.scala 43:79]
  wire  dontForward1 = _T & _T_1; // @[ISU.scala 43:57]
  wire  _T_2 = io_in_0_bits_ctrl_rfSrc1 != 5'h0; // @[ISU.scala 40:69]
  wire  _T_3 = io_in_0_bits_ctrl_rfSrc1 == io_forward_wb_rfDest; // @[ISU.scala 40:88]
  wire  _T_4 = _T_2 & _T_3; // @[ISU.scala 40:78]
  wire  src1DependEX = _T_4 & forwardRfWen; // @[ISU.scala 40:100]
  wire  _T_5 = io_in_0_bits_ctrl_rfSrc2 != 5'h0; // @[ISU.scala 40:69]
  wire  _T_6 = io_in_0_bits_ctrl_rfSrc2 == io_forward_wb_rfDest; // @[ISU.scala 40:88]
  wire  _T_7 = _T_5 & _T_6; // @[ISU.scala 40:78]
  wire  src2DependEX = _T_7 & forwardRfWen; // @[ISU.scala 40:100]
  wire  _T_9 = io_in_0_bits_ctrl_rfSrc1 == io_wb_rfDest; // @[ISU.scala 40:88]
  wire  _T_10 = _T_2 & _T_9; // @[ISU.scala 40:78]
  wire  src1DependWB = _T_10 & io_wb_rfWen; // @[ISU.scala 40:100]
  wire  _T_12 = io_in_0_bits_ctrl_rfSrc2 == io_wb_rfDest; // @[ISU.scala 40:88]
  wire  _T_13 = _T_5 & _T_12; // @[ISU.scala 40:78]
  wire  src2DependWB = _T_13 & io_wb_rfWen; // @[ISU.scala 40:100]
  wire  _T_14 = ~dontForward1; // @[ISU.scala 49:46]
  wire  src1ForwardNextCycle = src1DependEX & _T_14; // @[ISU.scala 49:43]
  wire  src2ForwardNextCycle = src2DependEX & _T_14; // @[ISU.scala 50:43]
  wire  _T_16 = ~src1DependEX; // @[ISU.scala 51:55]
  wire  _T_17 = dontForward1 ? _T_16 : 1'h1; // @[ISU.scala 51:40]
  wire  src1Forward = src1DependWB & _T_17; // @[ISU.scala 51:34]
  wire  _T_18 = ~src2DependEX; // @[ISU.scala 52:55]
  wire  _T_19 = dontForward1 ? _T_18 : 1'h1; // @[ISU.scala 52:40]
  wire  src2Forward = src2DependWB & _T_19; // @[ISU.scala 52:34]
  reg [31:0] _T_20; // @[RF.scala 36:21]
  wire [31:0] _T_21 = _T_20 >> io_in_0_bits_ctrl_rfSrc1; // @[RF.scala 37:37]
  wire  _T_23 = ~_T_21[0]; // @[ISU.scala 55:19]
  wire  _T_24 = _T_23 | src1ForwardNextCycle; // @[ISU.scala 55:38]
  wire  src1Ready = _T_24 | src1Forward; // @[ISU.scala 55:62]
  wire [31:0] _T_25 = _T_20 >> io_in_0_bits_ctrl_rfSrc2; // @[RF.scala 37:37]
  wire  _T_27 = ~_T_25[0]; // @[ISU.scala 56:19]
  wire  _T_28 = _T_27 | src2ForwardNextCycle; // @[ISU.scala 56:38]
  wire  src2Ready = _T_28 | src2Forward; // @[ISU.scala 56:62]
  wire  _T_29 = io_in_0_valid & src1Ready; // @[ISU.scala 57:34]
  wire [24:0] _T_35 = io_in_0_bits_cf_pc[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_36 = {_T_35,io_in_0_bits_cf_pc}; // @[Cat.scala 29:58]
  wire  _T_37 = ~src1ForwardNextCycle; // @[ISU.scala 65:21]
  wire  _T_38 = src1Forward & _T_37; // @[ISU.scala 65:18]
  wire  _T_39 = ~io_in_0_bits_ctrl_src1Type; // @[ISU.scala 66:35]
  wire  _T_41 = _T_39 & _T_37; // @[ISU.scala 66:51]
  wire  _T_42 = ~src1Forward; // @[ISU.scala 66:79]
  wire  _T_43 = _T_41 & _T_42; // @[ISU.scala 66:76]
  wire  _T_44 = io_in_0_bits_ctrl_rfSrc1 == 5'h0; // @[RF.scala 31:42]
  wire [63:0] _T_46 = _T_44 ? 64'h0 : _T_31__T_45_data; // @[RF.scala 31:36]
  wire [63:0] _T_47 = io_in_0_bits_ctrl_src1Type ? _T_36 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_48 = src1ForwardNextCycle ? io_forward_wb_rfData : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_49 = _T_38 ? io_wb_rfData : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_50 = _T_43 ? _T_46 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_51 = _T_47 | _T_48; // @[Mux.scala 27:72]
  wire [63:0] _T_52 = _T_51 | _T_49; // @[Mux.scala 27:72]
  wire  _T_56 = ~src2ForwardNextCycle; // @[ISU.scala 71:21]
  wire  _T_57 = src2Forward & _T_56; // @[ISU.scala 71:18]
  wire  _T_58 = ~io_in_0_bits_ctrl_src2Type; // @[ISU.scala 72:35]
  wire  _T_60 = _T_58 & _T_56; // @[ISU.scala 72:52]
  wire  _T_61 = ~src2Forward; // @[ISU.scala 72:80]
  wire  _T_62 = _T_60 & _T_61; // @[ISU.scala 72:77]
  wire  _T_63 = io_in_0_bits_ctrl_rfSrc2 == 5'h0; // @[RF.scala 31:42]
  wire [63:0] _T_65 = _T_63 ? 64'h0 : _T_31__T_64_data; // @[RF.scala 31:36]
  wire [63:0] _T_66 = io_in_0_bits_ctrl_src2Type ? io_in_0_bits_data_imm : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_67 = src2ForwardNextCycle ? io_forward_wb_rfData : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_68 = _T_57 ? io_wb_rfData : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_69 = _T_62 ? _T_65 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_70 = _T_66 | _T_67; // @[Mux.scala 27:72]
  wire [63:0] _T_71 = _T_70 | _T_68; // @[Mux.scala 27:72]
  wire  _T_76 = io_wb_rfDest != 5'h0; // @[ISU.scala 40:69]
  wire  _T_77 = io_wb_rfDest == io_forward_wb_rfDest; // @[ISU.scala 40:88]
  wire  _T_78 = _T_76 & _T_77; // @[ISU.scala 40:78]
  wire  _T_79 = _T_78 & forwardRfWen; // @[ISU.scala 40:100]
  wire  _T_80 = ~_T_79; // @[ISU.scala 84:40]
  wire  _T_81 = io_wb_rfWen & _T_80; // @[ISU.scala 84:37]
  wire [62:0] _T_82 = 63'h1 << io_wb_rfDest; // @[RF.scala 38:39]
  wire [31:0] wbClearMask = _T_81 ? _T_82[31:0] : 32'h0; // @[ISU.scala 84:24]
  wire  _T_84 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire [62:0] _T_85 = 63'h1 << io_in_0_bits_ctrl_rfDest; // @[RF.scala 38:39]
  wire [31:0] isuFireSetMask = _T_84 ? _T_85[31:0] : 32'h0; // @[ISU.scala 86:27]
  wire [31:0] _T_93 = ~wbClearMask; // @[RF.scala 44:26]
  wire [31:0] _T_94 = _T_20 & _T_93; // @[RF.scala 44:24]
  wire [31:0] _T_95 = _T_94 | isuFireSetMask; // @[RF.scala 44:38]
  wire [31:0] _T_97 = {_T_95[31:1],1'h0}; // @[Cat.scala 29:58]
  wire  _T_98 = ~io_in_0_valid; // @[ISU.scala 90:21]
  wire  _T_111 = ~io_out_valid; // @[ISU.scala 96:43]
  wire  _T_112 = io_in_0_valid & _T_111; // @[ISU.scala 96:40]
  wire  _T_114 = ~_T_84; // @[ISU.scala 97:41]
  wire  _T_115 = io_out_valid & _T_114; // @[ISU.scala 97:38]
  wire  _T_116 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign _T_31__T_45_addr = io_in_0_bits_ctrl_rfSrc1;
  assign _T_31__T_45_data = _T_31[_T_31__T_45_addr]; // @[RF.scala 30:15]
  assign _T_31__T_64_addr = io_in_0_bits_ctrl_rfSrc2;
  assign _T_31__T_64_data = _T_31[_T_31__T_64_addr]; // @[RF.scala 30:15]
  assign _T_31__T_74_data = io_wb_rfData;
  assign _T_31__T_74_addr = io_wb_rfDest;
  assign _T_31__T_74_mask = 1'h1;
  assign _T_31__T_74_en = io_wb_rfWen;
  assign io_in_0_ready = _T_98 | _T_84; // @[ISU.scala 90:18]
  assign io_out_valid = _T_29 & src2Ready; // @[ISU.scala 57:16]
  assign io_out_bits_cf_instr = io_in_0_bits_cf_instr; // @[ISU.scala 76:18]
  assign io_out_bits_cf_pc = io_in_0_bits_cf_pc; // @[ISU.scala 76:18]
  assign io_out_bits_cf_pnpc = io_in_0_bits_cf_pnpc; // @[ISU.scala 76:18]
  assign io_out_bits_cf_exceptionVec_1 = io_in_0_bits_cf_exceptionVec_1; // @[ISU.scala 76:18]
  assign io_out_bits_cf_exceptionVec_2 = io_in_0_bits_cf_exceptionVec_2; // @[ISU.scala 76:18]
  assign io_out_bits_cf_exceptionVec_12 = io_in_0_bits_cf_exceptionVec_12; // @[ISU.scala 76:18]
  assign io_out_bits_cf_intrVec_0 = io_in_0_bits_cf_intrVec_0; // @[ISU.scala 76:18]
  assign io_out_bits_cf_intrVec_1 = io_in_0_bits_cf_intrVec_1; // @[ISU.scala 76:18]
  assign io_out_bits_cf_intrVec_2 = io_in_0_bits_cf_intrVec_2; // @[ISU.scala 76:18]
  assign io_out_bits_cf_intrVec_3 = io_in_0_bits_cf_intrVec_3; // @[ISU.scala 76:18]
  assign io_out_bits_cf_intrVec_4 = io_in_0_bits_cf_intrVec_4; // @[ISU.scala 76:18]
  assign io_out_bits_cf_intrVec_5 = io_in_0_bits_cf_intrVec_5; // @[ISU.scala 76:18]
  assign io_out_bits_cf_intrVec_6 = io_in_0_bits_cf_intrVec_6; // @[ISU.scala 76:18]
  assign io_out_bits_cf_intrVec_7 = io_in_0_bits_cf_intrVec_7; // @[ISU.scala 76:18]
  assign io_out_bits_cf_intrVec_8 = io_in_0_bits_cf_intrVec_8; // @[ISU.scala 76:18]
  assign io_out_bits_cf_intrVec_9 = io_in_0_bits_cf_intrVec_9; // @[ISU.scala 76:18]
  assign io_out_bits_cf_intrVec_10 = io_in_0_bits_cf_intrVec_10; // @[ISU.scala 76:18]
  assign io_out_bits_cf_intrVec_11 = io_in_0_bits_cf_intrVec_11; // @[ISU.scala 76:18]
  assign io_out_bits_cf_brIdx = io_in_0_bits_cf_brIdx; // @[ISU.scala 76:18]
  assign io_out_bits_cf_crossPageIPFFix = io_in_0_bits_cf_crossPageIPFFix; // @[ISU.scala 76:18]
  assign io_out_bits_ctrl_fuType = io_in_0_bits_ctrl_fuType; // @[ISU.scala 77:20]
  assign io_out_bits_ctrl_fuOpType = io_in_0_bits_ctrl_fuOpType; // @[ISU.scala 77:20]
  assign io_out_bits_ctrl_rfWen = io_in_0_bits_ctrl_rfWen; // @[ISU.scala 77:20]
  assign io_out_bits_ctrl_rfDest = io_in_0_bits_ctrl_rfDest; // @[ISU.scala 77:20]
  assign io_out_bits_data_src1 = _T_52 | _T_50; // @[ISU.scala 62:25]
  assign io_out_bits_data_src2 = _T_71 | _T_69; // @[ISU.scala 68:25]
  assign io_out_bits_data_imm = io_in_0_bits_data_imm; // @[ISU.scala 74:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {2{`RANDOM}};
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    _T_31[initvar] = _RAND_0[63:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_20 = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_31__T_74_en & _T_31__T_74_mask) begin
      _T_31[_T_31__T_74_addr] <= _T_31__T_74_data; // @[RF.scala 30:15]
    end
    if (reset) begin
      _T_20 <= 32'h0;
    end else if (io_flush) begin
      _T_20 <= 32'h0;
    end else begin
      _T_20 <= _T_97;
    end
  end
endmodule
module ALU(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [63:0] io_in_bits_src1,
  input  [63:0] io_in_bits_src2,
  input  [6:0]  io_in_bits_func,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits,
  input  [63:0] io_cfIn_instr,
  input  [38:0] io_cfIn_pc,
  input  [38:0] io_cfIn_pnpc,
  input  [3:0]  io_cfIn_brIdx,
  output [38:0] io_redirect_target,
  output        io_redirect_valid,
  input  [63:0] io_offset,
  output        _T_243_0_valid,
  output [38:0] _T_243_0_pc,
  output        _T_243_0_isMissPredict,
  output [38:0] _T_243_0_actualTarget,
  output        _T_243_0_actualTaken,
  output [6:0]  _T_243_0_fuOpType,
  output [1:0]  _T_243_0_btbType,
  output        _T_243_0_isRVC
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire  isAdderSub = ~io_in_bits_func[6]; // @[ALU.scala 86:20]
  wire [63:0] _T_2 = isAdderSub ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_3 = io_in_bits_src2 ^ _T_2; // @[ALU.scala 87:33]
  wire [64:0] _T_4 = io_in_bits_src1 + _T_3; // @[ALU.scala 87:24]
  wire [64:0] _GEN_0 = {{64'd0}, isAdderSub}; // @[ALU.scala 87:60]
  wire [64:0] adderRes = _T_4 + _GEN_0; // @[ALU.scala 87:60]
  wire [63:0] xorRes = io_in_bits_src1 ^ io_in_bits_src2; // @[ALU.scala 88:21]
  wire  sltu = ~adderRes[64]; // @[ALU.scala 89:14]
  wire  slt = xorRes[63] ^ sltu; // @[ALU.scala 90:28]
  wire [63:0] _T_10 = {32'h0,io_in_bits_src1[31:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_14 = io_in_bits_src1[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_15 = {_T_14,io_in_bits_src1[31:0]}; // @[Cat.scala 29:58]
  wire  _T_16 = 7'h25 == io_in_bits_func; // @[Mux.scala 80:60]
  wire [63:0] _T_17 = _T_16 ? _T_10 : io_in_bits_src1; // @[Mux.scala 80:57]
  wire  _T_18 = 7'h2d == io_in_bits_func; // @[Mux.scala 80:60]
  wire [63:0] shsrc1 = _T_18 ? _T_15 : _T_17; // @[Mux.scala 80:57]
  wire [5:0] shamt = io_in_bits_func[5] ? {{1'd0}, io_in_bits_src2[4:0]} : io_in_bits_src2[5:0]; // @[ALU.scala 96:18]
  wire [126:0] _GEN_1 = {{63'd0}, shsrc1}; // @[ALU.scala 98:33]
  wire [126:0] _T_23 = _GEN_1 << shamt; // @[ALU.scala 98:33]
  wire [63:0] _T_25 = {63'h0,slt}; // @[Cat.scala 29:58]
  wire [63:0] _T_26 = {63'h0,sltu}; // @[Cat.scala 29:58]
  wire [63:0] _T_27 = shsrc1 >> shamt; // @[ALU.scala 102:32]
  wire [63:0] _T_28 = io_in_bits_src1 | io_in_bits_src2; // @[ALU.scala 103:30]
  wire [63:0] _T_29 = io_in_bits_src1 & io_in_bits_src2; // @[ALU.scala 104:30]
  wire [63:0] _T_30 = _T_18 ? _T_15 : _T_17; // @[ALU.scala 105:32]
  wire [63:0] _T_32 = $signed(_T_30) >>> shamt; // @[ALU.scala 105:49]
  wire  _T_33 = 4'h1 == io_in_bits_func[3:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_34 = _T_33 ? {{1'd0}, _T_23[63:0]} : adderRes; // @[Mux.scala 80:57]
  wire  _T_35 = 4'h2 == io_in_bits_func[3:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_36 = _T_35 ? {{1'd0}, _T_25} : _T_34; // @[Mux.scala 80:57]
  wire  _T_37 = 4'h3 == io_in_bits_func[3:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_38 = _T_37 ? {{1'd0}, _T_26} : _T_36; // @[Mux.scala 80:57]
  wire  _T_39 = 4'h4 == io_in_bits_func[3:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_40 = _T_39 ? {{1'd0}, xorRes} : _T_38; // @[Mux.scala 80:57]
  wire  _T_41 = 4'h5 == io_in_bits_func[3:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_42 = _T_41 ? {{1'd0}, _T_27} : _T_40; // @[Mux.scala 80:57]
  wire  _T_43 = 4'h6 == io_in_bits_func[3:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_44 = _T_43 ? {{1'd0}, _T_28} : _T_42; // @[Mux.scala 80:57]
  wire  _T_45 = 4'h7 == io_in_bits_func[3:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_46 = _T_45 ? {{1'd0}, _T_29} : _T_44; // @[Mux.scala 80:57]
  wire  _T_47 = 4'hd == io_in_bits_func[3:0]; // @[Mux.scala 80:60]
  wire [64:0] res = _T_47 ? {{1'd0}, _T_32} : _T_46; // @[Mux.scala 80:57]
  wire [31:0] _T_52 = res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_53 = {_T_52,res[31:0]}; // @[Cat.scala 29:58]
  wire [64:0] aluRes = io_in_bits_func[5] ? {{1'd0}, _T_53} : res; // @[ALU.scala 107:19]
  wire  _T_54 = |xorRes; // @[ALU.scala 110:56]
  wire  _T_55 = ~_T_54; // @[ALU.scala 110:48]
  wire  isBranch = ~io_in_bits_func[3]; // @[ALU.scala 62:30]
  wire  isBru = io_in_bits_func[4]; // @[ALU.scala 61:31]
  wire  _T_58 = 2'h0 == io_in_bits_func[2:1]; // @[LookupTree.scala 24:34]
  wire  _T_59 = 2'h2 == io_in_bits_func[2:1]; // @[LookupTree.scala 24:34]
  wire  _T_60 = 2'h3 == io_in_bits_func[2:1]; // @[LookupTree.scala 24:34]
  wire  _T_61 = _T_58 & _T_55; // @[Mux.scala 27:72]
  wire  _T_62 = _T_59 & slt; // @[Mux.scala 27:72]
  wire  _T_63 = _T_60 & sltu; // @[Mux.scala 27:72]
  wire  _T_64 = _T_61 | _T_62; // @[Mux.scala 27:72]
  wire  _T_65 = _T_64 | _T_63; // @[Mux.scala 27:72]
  wire  taken = _T_65 ^ io_in_bits_func[0]; // @[ALU.scala 117:72]
  wire [63:0] _GEN_2 = {{25'd0}, io_cfIn_pc}; // @[ALU.scala 118:41]
  wire [63:0] _T_69 = _GEN_2 + io_offset; // @[ALU.scala 118:41]
  wire [64:0] _T_70 = isBranch ? {{1'd0}, _T_69} : adderRes; // @[ALU.scala 118:19]
  wire [38:0] target = _T_70[38:0]; // @[ALU.scala 118:63]
  wire  _T_71 = ~taken; // @[ALU.scala 119:26]
  wire  _T_72 = _T_71 & isBranch; // @[ALU.scala 119:33]
  wire  _T_75 = ~io_cfIn_brIdx[0]; // @[ALU.scala 119:64]
  wire  _T_76 = io_redirect_target != io_cfIn_pnpc; // @[ALU.scala 119:105]
  wire  _T_77 = _T_75 | _T_76; // @[ALU.scala 119:82]
  wire  predictWrong = _T_72 ? io_cfIn_brIdx[0] : _T_77; // @[ALU.scala 119:25]
  wire  isRVC = io_cfIn_instr[1:0] != 2'h3; // @[ALU.scala 120:35]
  wire  _T_80 = io_cfIn_instr[1:0] == 2'h3; // @[ALU.scala 121:29]
  wire  _T_81 = _T_80 | isRVC; // @[ALU.scala 121:41]
  wire  _T_82 = ~io_in_valid; // @[ALU.scala 121:53]
  wire  _T_83 = _T_81 | _T_82; // @[ALU.scala 121:50]
  wire  _T_85 = _T_83 | reset; // @[ALU.scala 121:9]
  wire  _T_86 = ~_T_85; // @[ALU.scala 121:9]
  wire  _T_89 = ~isRVC; // @[ALU.scala 122:55]
  wire [38:0] _T_104 = io_cfIn_pc + 39'h2; // @[ALU.scala 123:71]
  wire [38:0] _T_106 = io_cfIn_pc + 39'h4; // @[ALU.scala 123:89]
  wire [38:0] _T_107 = isRVC ? _T_104 : _T_106; // @[ALU.scala 123:52]
  wire  _T_109 = io_in_valid & isBru; // @[ALU.scala 125:30]
  wire  _T_110 = _T_109 & predictWrong; // @[ALU.scala 125:39]
  wire [24:0] _T_114 = io_cfIn_pc[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_115 = {_T_114,io_cfIn_pc}; // @[Cat.scala 29:58]
  wire [63:0] _T_117 = _T_115 + 64'h4; // @[ALU.scala 131:71]
  wire [63:0] _T_123 = _T_115 + 64'h2; // @[ALU.scala 131:108]
  wire [63:0] _T_124 = _T_89 ? _T_117 : _T_123; // @[ALU.scala 131:32]
  wire [64:0] _T_125 = isBru ? {{1'd0}, _T_124} : aluRes; // @[ALU.scala 131:21]
  wire  _T_147 = io_in_bits_func == 7'h58; // @[ALU.scala 135:162]
  wire  _T_148 = io_in_bits_func == 7'h5c; // @[ALU.scala 135:188]
  wire  _T_149 = _T_147 | _T_148; // @[ALU.scala 135:180]
  wire  _T_150 = io_in_bits_func == 7'h5a; // @[ALU.scala 135:214]
  wire  _T_151 = io_in_bits_func == 7'h5e; // @[ALU.scala 135:239]
  wire  _T_178 = 7'h5c == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_179 = 7'h5e == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_180 = 7'h58 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_181 = 7'h5a == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire [1:0] _T_189 = _T_179 ? 2'h3 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _T_191 = _T_181 ? 2'h2 : 2'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_3 = {{1'd0}, _T_178}; // @[Mux.scala 27:72]
  wire [1:0] _T_198 = _GEN_3 | _T_189; // @[Mux.scala 27:72]
  wire [1:0] _GEN_4 = {{1'd0}, _T_180}; // @[Mux.scala 27:72]
  wire [1:0] _T_199 = _T_198 | _GEN_4; // @[Mux.scala 27:72]
  reg  _T_243_valid; // @[ALU.scala 158:34]
  reg [38:0] _T_243_pc; // @[ALU.scala 158:34]
  reg  _T_243_isMissPredict; // @[ALU.scala 158:34]
  reg [38:0] _T_243_actualTarget; // @[ALU.scala 158:34]
  reg  _T_243_actualTaken; // @[ALU.scala 158:34]
  reg [6:0] _T_243_fuOpType; // @[ALU.scala 158:34]
  reg [1:0] _T_243_btbType; // @[ALU.scala 158:34]
  reg  _T_243_isRVC; // @[ALU.scala 158:34]
  wire  _T_245 = ~predictWrong; // @[ALU.scala 160:35]
  wire  _T_246 = _T_109 & _T_245; // @[ALU.scala 160:32]
  wire  _T_249 = _T_246 & isBranch; // @[ALU.scala 162:33]
  wire  _T_250 = _T_110 & isBranch; // @[ALU.scala 163:33]
  wire  _T_253 = io_cfIn_pc[2:0] == 3'h0; // @[ALU.scala 164:63]
  wire  _T_254 = _T_250 & _T_253; // @[ALU.scala 164:45]
  wire  _T_255 = _T_254 & isRVC; // @[ALU.scala 164:73]
  wire  _T_261 = _T_254 & _T_89; // @[ALU.scala 165:73]
  wire  _T_264 = io_cfIn_pc[2:0] == 3'h2; // @[ALU.scala 166:63]
  wire  _T_265 = _T_250 & _T_264; // @[ALU.scala 166:45]
  wire  _T_266 = _T_265 & isRVC; // @[ALU.scala 166:73]
  wire  _T_272 = _T_265 & _T_89; // @[ALU.scala 167:73]
  wire  _T_275 = io_cfIn_pc[2:0] == 3'h4; // @[ALU.scala 168:63]
  wire  _T_276 = _T_250 & _T_275; // @[ALU.scala 168:45]
  wire  _T_277 = _T_276 & isRVC; // @[ALU.scala 168:73]
  wire  _T_283 = _T_276 & _T_89; // @[ALU.scala 169:73]
  wire  _T_286 = io_cfIn_pc[2:0] == 3'h6; // @[ALU.scala 170:63]
  wire  _T_287 = _T_250 & _T_286; // @[ALU.scala 170:45]
  wire  _T_288 = _T_287 & isRVC; // @[ALU.scala 170:73]
  wire  _T_294 = _T_287 & _T_89; // @[ALU.scala 171:73]
  wire  _T_298 = _T_246 & _T_149; // @[ALU.scala 172:33]
  wire  _T_302 = _T_110 & _T_149; // @[ALU.scala 173:33]
  wire  _T_304 = _T_246 & _T_150; // @[ALU.scala 174:33]
  wire  _T_306 = _T_110 & _T_150; // @[ALU.scala 175:33]
  wire  _T_308 = _T_246 & _T_151; // @[ALU.scala 176:33]
  wire  _T_310 = _T_110 & _T_151; // @[ALU.scala 177:33]
  assign io_out_valid = io_in_valid; // @[ALU.scala 145:16]
  assign io_out_bits = _T_125[63:0]; // @[ALU.scala 131:15]
  assign io_redirect_target = _T_72 ? _T_107 : target; // @[ALU.scala 123:22]
  assign io_redirect_valid = _T_109 & predictWrong; // @[ALU.scala 125:21]
  assign _T_243_0_valid = _T_243_valid;
  assign _T_243_0_pc = _T_243_pc;
  assign _T_243_0_isMissPredict = _T_243_isMissPredict;
  assign _T_243_0_actualTarget = _T_243_actualTarget;
  assign _T_243_0_actualTaken = _T_243_actualTaken;
  assign _T_243_0_fuOpType = _T_243_fuOpType;
  assign _T_243_0_btbType = _T_243_btbType;
  assign _T_243_0_isRVC = _T_243_isRVC;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_243_valid = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  _T_243_pc = _RAND_1[38:0];
  _RAND_2 = {1{`RANDOM}};
  _T_243_isMissPredict = _RAND_2[0:0];
  _RAND_3 = {2{`RANDOM}};
  _T_243_actualTarget = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  _T_243_actualTaken = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_243_fuOpType = _RAND_5[6:0];
  _RAND_6 = {1{`RANDOM}};
  _T_243_btbType = _RAND_6[1:0];
  _RAND_7 = {1{`RANDOM}};
  _T_243_isRVC = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_243_valid <= io_in_valid & isBru;
    _T_243_pc <= io_cfIn_pc;
    if (_T_72) begin
      _T_243_isMissPredict <= io_cfIn_brIdx[0];
    end else begin
      _T_243_isMissPredict <= _T_77;
    end
    _T_243_actualTarget <= _T_70[38:0];
    _T_243_actualTaken <= _T_65 ^ io_in_bits_func[0];
    _T_243_fuOpType <= io_in_bits_func;
    _T_243_btbType <= _T_199 | _T_191;
    _T_243_isRVC <= io_cfIn_instr[1:0] != 2'h3;
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_86) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ALU.scala:121 assert(io.cfIn.instr(1,0) === \"b11\".U || isRVC || !valid)\n"); // @[ALU.scala 121:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_86) begin
          $fatal; // @[ALU.scala 121:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module LSExecUnit(
  input         clock,
  input         reset,
  input         io__in_valid,
  input  [63:0] io__in_bits_src1,
  input  [6:0]  io__in_bits_func,
  input         io__out_ready,
  output        io__out_valid,
  output [63:0] io__out_bits,
  input  [63:0] io__wdata,
  input         io__dmem_req_ready,
  output        io__dmem_req_valid,
  output [38:0] io__dmem_req_bits_addr,
  output [2:0]  io__dmem_req_bits_size,
  output [3:0]  io__dmem_req_bits_cmd,
  output [7:0]  io__dmem_req_bits_wmask,
  output [63:0] io__dmem_req_bits_wdata,
  output        io__dmem_resp_ready,
  input         io__dmem_resp_valid,
  input  [63:0] io__dmem_resp_bits_rdata,
  output        io__isMMIO,
  output        io__dtlbPF,
  output        io__loadAddrMisaligned,
  output        io__storeAddrMisaligned,
  input         DTLBPF,
  input         DTLBENABLE,
  input         ISAMO2,
  output [63:0] io_in_bits_src1,
  input         DTLBFINISH
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] addrLatch; // @[UnpipelinedLSU.scala 333:26]
  wire  isStore = io__in_valid & io__in_bits_func[3]; // @[UnpipelinedLSU.scala 334:23]
  wire  _T_1 = ~isStore; // @[UnpipelinedLSU.scala 335:21]
  wire  _T_2 = io__in_bits_func != 7'h3; // @[UnpipelinedLSU.scala 335:39]
  wire  partialLoad = _T_1 & _T_2; // @[UnpipelinedLSU.scala 335:30]
  reg [1:0] state; // @[UnpipelinedLSU.scala 338:22]
  wire  _T_3 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_4 = io__dmem_req_ready & io__dmem_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_5 = _T_4 & DTLBENABLE; // @[UnpipelinedLSU.scala 353:29]
  wire  _T_7 = ~DTLBENABLE; // @[UnpipelinedLSU.scala 354:32]
  wire  _T_8 = _T_4 & _T_7; // @[UnpipelinedLSU.scala 354:29]
  wire  _T_9 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_10 = DTLBFINISH & DTLBPF; // @[UnpipelinedLSU.scala 358:24]
  wire  _T_11 = ~DTLBPF; // @[UnpipelinedLSU.scala 359:27]
  wire  _T_12 = DTLBFINISH & _T_11; // @[UnpipelinedLSU.scala 359:24]
  wire  _T_13 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_14 = io__dmem_resp_ready & io__dmem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_16 = 2'h3 == state; // @[Conditional.scala 37:30]
  wire [63:0] _T_55 = {io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0],io__wdata[7:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_58 = {io__wdata[15:0],io__wdata[15:0],io__wdata[15:0],io__wdata[15:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_60 = {io__wdata[31:0],io__wdata[31:0]}; // @[Cat.scala 29:58]
  wire  _T_61 = 2'h0 == io__in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_62 = 2'h1 == io__in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_63 = 2'h2 == io__in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_64 = 2'h3 == io__in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire [63:0] _T_65 = _T_61 ? _T_55 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_66 = _T_62 ? _T_58 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_67 = _T_63 ? _T_60 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_68 = _T_64 ? io__wdata : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_69 = _T_65 | _T_66; // @[Mux.scala 27:72]
  wire [63:0] _T_70 = _T_69 | _T_67; // @[Mux.scala 27:72]
  wire [1:0] _T_77 = _T_62 ? 2'h3 : 2'h0; // @[Mux.scala 27:72]
  wire [3:0] _T_78 = _T_63 ? 4'hf : 4'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_79 = _T_64 ? 8'hff : 8'h0; // @[Mux.scala 27:72]
  wire [1:0] _GEN_13 = {{1'd0}, _T_61}; // @[Mux.scala 27:72]
  wire [1:0] _T_80 = _GEN_13 | _T_77; // @[Mux.scala 27:72]
  wire [3:0] _GEN_14 = {{2'd0}, _T_80}; // @[Mux.scala 27:72]
  wire [3:0] _T_81 = _GEN_14 | _T_78; // @[Mux.scala 27:72]
  wire [7:0] _GEN_15 = {{4'd0}, _T_81}; // @[Mux.scala 27:72]
  wire [7:0] _T_82 = _GEN_15 | _T_79; // @[Mux.scala 27:72]
  wire [14:0] _GEN_16 = {{7'd0}, _T_82}; // @[UnpipelinedLSU.scala 306:8]
  wire [14:0] reqWmask = _GEN_16 << io__in_bits_src1[2:0]; // @[UnpipelinedLSU.scala 306:8]
  wire  _T_86 = state == 2'h0; // @[UnpipelinedLSU.scala 379:37]
  wire  _T_87 = io__in_valid & _T_86; // @[UnpipelinedLSU.scala 379:27]
  wire  _T_88 = ~io__loadAddrMisaligned; // @[UnpipelinedLSU.scala 379:52]
  wire  _T_89 = _T_87 & _T_88; // @[UnpipelinedLSU.scala 379:49]
  wire  _T_90 = ~io__storeAddrMisaligned; // @[UnpipelinedLSU.scala 379:78]
  wire  _T_92 = state != 2'h0; // @[UnpipelinedLSU.scala 382:40]
  wire  _T_93 = DTLBPF & _T_92; // @[UnpipelinedLSU.scala 382:31]
  wire  _T_94 = _T_93 | io__loadAddrMisaligned; // @[UnpipelinedLSU.scala 382:51]
  wire  _T_95 = _T_94 | io__storeAddrMisaligned; // @[UnpipelinedLSU.scala 382:76]
  wire  _T_96 = state == 2'h3; // @[UnpipelinedLSU.scala 382:134]
  wire  _T_98 = state == 2'h2; // @[UnpipelinedLSU.scala 382:180]
  wire  _T_99 = _T_14 & _T_98; // @[UnpipelinedLSU.scala 382:170]
  wire  _T_100 = partialLoad ? _T_96 : _T_99; // @[UnpipelinedLSU.scala 382:114]
  reg [63:0] rdataLatch; // @[UnpipelinedLSU.scala 388:27]
  wire  _T_124 = 3'h0 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_125 = 3'h1 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_126 = 3'h2 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_127 = 3'h3 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_128 = 3'h4 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_129 = 3'h5 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_130 = 3'h6 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire  _T_131 = 3'h7 == addrLatch[2:0]; // @[LookupTree.scala 24:34]
  wire [63:0] _T_132 = _T_124 ? rdataLatch : 64'h0; // @[Mux.scala 27:72]
  wire [55:0] _T_133 = _T_125 ? rdataLatch[63:8] : 56'h0; // @[Mux.scala 27:72]
  wire [47:0] _T_134 = _T_126 ? rdataLatch[63:16] : 48'h0; // @[Mux.scala 27:72]
  wire [39:0] _T_135 = _T_127 ? rdataLatch[63:24] : 40'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_136 = _T_128 ? rdataLatch[63:32] : 32'h0; // @[Mux.scala 27:72]
  wire [23:0] _T_137 = _T_129 ? rdataLatch[63:40] : 24'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_138 = _T_130 ? rdataLatch[63:48] : 16'h0; // @[Mux.scala 27:72]
  wire [7:0] _T_139 = _T_131 ? rdataLatch[63:56] : 8'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_17 = {{8'd0}, _T_133}; // @[Mux.scala 27:72]
  wire [63:0] _T_140 = _T_132 | _GEN_17; // @[Mux.scala 27:72]
  wire [63:0] _GEN_18 = {{16'd0}, _T_134}; // @[Mux.scala 27:72]
  wire [63:0] _T_141 = _T_140 | _GEN_18; // @[Mux.scala 27:72]
  wire [63:0] _GEN_19 = {{24'd0}, _T_135}; // @[Mux.scala 27:72]
  wire [63:0] _T_142 = _T_141 | _GEN_19; // @[Mux.scala 27:72]
  wire [63:0] _GEN_20 = {{32'd0}, _T_136}; // @[Mux.scala 27:72]
  wire [63:0] _T_143 = _T_142 | _GEN_20; // @[Mux.scala 27:72]
  wire [63:0] _GEN_21 = {{40'd0}, _T_137}; // @[Mux.scala 27:72]
  wire [63:0] _T_144 = _T_143 | _GEN_21; // @[Mux.scala 27:72]
  wire [63:0] _GEN_22 = {{48'd0}, _T_138}; // @[Mux.scala 27:72]
  wire [63:0] _T_145 = _T_144 | _GEN_22; // @[Mux.scala 27:72]
  wire [63:0] _GEN_23 = {{56'd0}, _T_139}; // @[Mux.scala 27:72]
  wire [63:0] rdataSel = _T_145 | _GEN_23; // @[Mux.scala 27:72]
  wire [55:0] _T_166 = rdataSel[7] ? 56'hffffffffffffff : 56'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_167 = {_T_166,rdataSel[7:0]}; // @[Cat.scala 29:58]
  wire [47:0] _T_171 = rdataSel[15] ? 48'hffffffffffff : 48'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_172 = {_T_171,rdataSel[15:0]}; // @[Cat.scala 29:58]
  wire [31:0] _T_176 = rdataSel[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_177 = {_T_176,rdataSel[31:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_179 = {56'h0,rdataSel[7:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_181 = {48'h0,rdataSel[15:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_183 = {32'h0,rdataSel[31:0]}; // @[Cat.scala 29:58]
  wire  _T_184 = 7'h0 == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_185 = 7'h1 == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_186 = 7'h2 == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_187 = 7'h4 == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_188 = 7'h5 == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_189 = 7'h6 == io__in_bits_func; // @[LookupTree.scala 24:34]
  wire [63:0] _T_190 = _T_184 ? _T_167 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_191 = _T_185 ? _T_172 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_192 = _T_186 ? _T_177 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_193 = _T_187 ? _T_179 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_194 = _T_188 ? _T_181 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_195 = _T_189 ? _T_183 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_196 = _T_190 | _T_191; // @[Mux.scala 27:72]
  wire [63:0] _T_197 = _T_196 | _T_192; // @[Mux.scala 27:72]
  wire [63:0] _T_198 = _T_197 | _T_193; // @[Mux.scala 27:72]
  wire [63:0] _T_199 = _T_198 | _T_194; // @[Mux.scala 27:72]
  wire [63:0] rdataPartialLoad = _T_199 | _T_195; // @[Mux.scala 27:72]
  wire  _T_203 = ~io__in_bits_src1[0]; // @[UnpipelinedLSU.scala 416:27]
  wire  _T_205 = io__in_bits_src1[1:0] == 2'h0; // @[UnpipelinedLSU.scala 417:29]
  wire  _T_207 = io__in_bits_src1[2:0] == 3'h0; // @[UnpipelinedLSU.scala 418:29]
  wire  _T_213 = _T_62 & _T_203; // @[Mux.scala 27:72]
  wire  _T_214 = _T_63 & _T_205; // @[Mux.scala 27:72]
  wire  _T_215 = _T_64 & _T_207; // @[Mux.scala 27:72]
  wire  _T_216 = _T_61 | _T_213; // @[Mux.scala 27:72]
  wire  _T_217 = _T_216 | _T_214; // @[Mux.scala 27:72]
  wire  addrAligned = _T_217 | _T_215; // @[Mux.scala 27:72]
  wire  _T_222 = io__in_valid & _T_1; // @[UnpipelinedLSU.scala 429:35]
  wire  _T_223 = ~ISAMO2; // @[UnpipelinedLSU.scala 429:50]
  wire  _T_224 = _T_222 & _T_223; // @[UnpipelinedLSU.scala 429:47]
  wire  _T_225 = ~addrAligned; // @[UnpipelinedLSU.scala 429:60]
  wire  _T_227 = isStore | ISAMO2; // @[UnpipelinedLSU.scala 430:47]
  wire  _T_228 = io__in_valid & _T_227; // @[UnpipelinedLSU.scala 430:35]
  wire  _T_242 = ~io__dmem_req_bits_cmd[0]; // @[SimpleBus.scala 73:18]
  wire  _T_244 = ~io__dmem_req_bits_cmd[3]; // @[SimpleBus.scala 73:29]
  wire  _T_245 = _T_242 & _T_244; // @[SimpleBus.scala 73:26]
  wire  _T_246 = io__dmem_req_valid & _T_245; // @[SimpleBus.scala 104:29]
  wire  _T_248 = _T_246 & _T_4; // @[UnpipelinedLSU.scala 434:39]
  reg  _T_256; // @[StopWatch.scala 24:20]
  wire  _GEN_9 = _T_246 | _T_256; // @[StopWatch.scala 30:20]
  wire  _T_258 = io__dmem_req_valid & io__dmem_req_bits_cmd[0]; // @[SimpleBus.scala 103:29]
  reg  _T_260; // @[StopWatch.scala 24:20]
  wire  _GEN_11 = _T_258 | _T_260; // @[StopWatch.scala 30:20]
  assign io__out_valid = _T_95 | _T_100; // @[UnpipelinedLSU.scala 382:16]
  assign io__out_bits = partialLoad ? rdataPartialLoad : io__dmem_resp_bits_rdata; // @[UnpipelinedLSU.scala 421:15]
  assign io__dmem_req_valid = _T_89 & _T_90; // @[UnpipelinedLSU.scala 379:18]
  assign io__dmem_req_bits_addr = io__in_bits_src1[38:0]; // @[SimpleBus.scala 64:15]
  assign io__dmem_req_bits_size = {{1'd0}, io__in_bits_func[1:0]}; // @[SimpleBus.scala 66:15]
  assign io__dmem_req_bits_cmd = {{3'd0}, isStore}; // @[SimpleBus.scala 65:14]
  assign io__dmem_req_bits_wmask = reqWmask[7:0]; // @[SimpleBus.scala 68:16]
  assign io__dmem_req_bits_wdata = _T_70 | _T_68; // @[SimpleBus.scala 67:16]
  assign io__dmem_resp_ready = 1'h1; // @[UnpipelinedLSU.scala 380:19]
  assign io__isMMIO = 1'h0;
  assign io__dtlbPF = DTLBPF; // @[UnpipelinedLSU.scala 349:13]
  assign io__loadAddrMisaligned = _T_224 & _T_225; // @[UnpipelinedLSU.scala 429:25]
  assign io__storeAddrMisaligned = _T_228 & _T_225; // @[UnpipelinedLSU.scala 430:26]
  assign io_in_bits_src1 = io__in_bits_src1;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  addrLatch = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[1:0];
  _RAND_2 = {2{`RANDOM}};
  rdataLatch = _RAND_2[63:0];
  _RAND_3 = {1{`RANDOM}};
  _T_256 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_260 = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    addrLatch <= io__in_bits_src1;
    if (reset) begin
      state <= 2'h0;
    end else if (_T_3) begin
      if (_T_8) begin
        state <= 2'h2;
      end else if (_T_5) begin
        state <= 2'h1;
      end
    end else if (_T_9) begin
      if (_T_12) begin
        state <= 2'h2;
      end else if (_T_10) begin
        state <= 2'h0;
      end
    end else if (_T_13) begin
      if (_T_14) begin
        if (partialLoad) begin
          state <= 2'h3;
        end else begin
          state <= 2'h0;
        end
      end
    end else if (_T_16) begin
      state <= 2'h0;
    end
    rdataLatch <= io__dmem_resp_bits_rdata;
    if (reset) begin
      _T_256 <= 1'h0;
    end else if (_T_14) begin
      _T_256 <= 1'h0;
    end else begin
      _T_256 <= _GEN_9;
    end
    if (reset) begin
      _T_260 <= 1'h0;
    end else if (_T_14) begin
      _T_260 <= 1'h0;
    end else begin
      _T_260 <= _GEN_11;
    end
  end
endmodule
module AtomALU(
  input  [63:0] io_src1,
  input  [63:0] io_src2,
  input  [6:0]  io_func,
  input         io_isWordOp,
  output [63:0] io_result
);
  wire  isAdderSub = ~io_func[6]; // @[LSU.scala 184:20]
  wire [63:0] _T_2 = isAdderSub ? 64'hffffffffffffffff : 64'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_3 = io_src2 ^ _T_2; // @[LSU.scala 185:33]
  wire [64:0] _T_4 = io_src1 + _T_3; // @[LSU.scala 185:24]
  wire [64:0] _GEN_0 = {{64'd0}, isAdderSub}; // @[LSU.scala 185:60]
  wire [64:0] adderRes = _T_4 + _GEN_0; // @[LSU.scala 185:60]
  wire [63:0] xorRes = io_src1 ^ io_src2; // @[LSU.scala 186:21]
  wire  sltu = ~adderRes[64]; // @[LSU.scala 187:14]
  wire  slt = xorRes[63] ^ sltu; // @[LSU.scala 188:28]
  wire [63:0] _T_9 = io_src1 & io_src2; // @[LSU.scala 194:32]
  wire [63:0] _T_10 = io_src1 | io_src2; // @[LSU.scala 195:32]
  wire [63:0] _T_12 = slt ? io_src1 : io_src2; // @[LSU.scala 196:29]
  wire [63:0] _T_14 = slt ? io_src2 : io_src1; // @[LSU.scala 197:29]
  wire [63:0] _T_16 = sltu ? io_src1 : io_src2; // @[LSU.scala 198:29]
  wire [63:0] _T_18 = sltu ? io_src2 : io_src1; // @[LSU.scala 199:29]
  wire  _T_19 = 6'h22 == io_func[5:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_20 = _T_19 ? {{1'd0}, io_src2} : adderRes; // @[Mux.scala 80:57]
  wire  _T_21 = 6'h24 == io_func[5:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_22 = _T_21 ? {{1'd0}, xorRes} : _T_20; // @[Mux.scala 80:57]
  wire  _T_23 = 6'h25 == io_func[5:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_24 = _T_23 ? {{1'd0}, _T_9} : _T_22; // @[Mux.scala 80:57]
  wire  _T_25 = 6'h26 == io_func[5:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_26 = _T_25 ? {{1'd0}, _T_10} : _T_24; // @[Mux.scala 80:57]
  wire  _T_27 = 6'h37 == io_func[5:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_28 = _T_27 ? {{1'd0}, _T_12} : _T_26; // @[Mux.scala 80:57]
  wire  _T_29 = 6'h30 == io_func[5:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_30 = _T_29 ? {{1'd0}, _T_14} : _T_28; // @[Mux.scala 80:57]
  wire  _T_31 = 6'h31 == io_func[5:0]; // @[Mux.scala 80:60]
  wire [64:0] _T_32 = _T_31 ? {{1'd0}, _T_16} : _T_30; // @[Mux.scala 80:57]
  wire  _T_33 = 6'h32 == io_func[5:0]; // @[Mux.scala 80:60]
  wire [64:0] res = _T_33 ? {{1'd0}, _T_18} : _T_32; // @[Mux.scala 80:57]
  wire [31:0] _T_37 = res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_38 = {_T_37,res[31:0]}; // @[Cat.scala 29:58]
  assign io_result = io_isWordOp ? _T_38 : res[63:0]; // @[LSU.scala 202:13]
endmodule
module UnpipelinedLSU(
  input         clock,
  input         reset,
  input         io__in_valid,
  input  [63:0] io__in_bits_src1,
  input  [63:0] io__in_bits_src2,
  input  [6:0]  io__in_bits_func,
  input         io__out_ready,
  output        io__out_valid,
  output [63:0] io__out_bits,
  input  [63:0] io__wdata,
  input  [31:0] io__instr,
  input         io__dmem_req_ready,
  output        io__dmem_req_valid,
  output [38:0] io__dmem_req_bits_addr,
  output [2:0]  io__dmem_req_bits_size,
  output [3:0]  io__dmem_req_bits_cmd,
  output [7:0]  io__dmem_req_bits_wmask,
  output [63:0] io__dmem_req_bits_wdata,
  input         io__dmem_resp_valid,
  input  [63:0] io__dmem_resp_bits_rdata,
  output        io__dtlbPF,
  output        io__loadAddrMisaligned,
  output        io__storeAddrMisaligned,
  output        setLr_0,
  input         DTLBPF,
  output        amoReq_0,
  input         DTLBENABLE,
  output [63:0] io_in_bits_src1,
  input         DTLBFINISH,
  output [63:0] setLrAddr_0,
  output        setLrVal_0,
  input  [63:0] lr_addr
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  lsExecUnit_clock; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_reset; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__in_valid; // @[UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io__in_bits_src1; // @[UnpipelinedLSU.scala 47:28]
  wire [6:0] lsExecUnit_io__in_bits_func; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__out_ready; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__out_valid; // @[UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io__out_bits; // @[UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io__wdata; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__dmem_req_ready; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__dmem_req_valid; // @[UnpipelinedLSU.scala 47:28]
  wire [38:0] lsExecUnit_io__dmem_req_bits_addr; // @[UnpipelinedLSU.scala 47:28]
  wire [2:0] lsExecUnit_io__dmem_req_bits_size; // @[UnpipelinedLSU.scala 47:28]
  wire [3:0] lsExecUnit_io__dmem_req_bits_cmd; // @[UnpipelinedLSU.scala 47:28]
  wire [7:0] lsExecUnit_io__dmem_req_bits_wmask; // @[UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io__dmem_req_bits_wdata; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__dmem_resp_ready; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__dmem_resp_valid; // @[UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io__dmem_resp_bits_rdata; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__isMMIO; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__dtlbPF; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__loadAddrMisaligned; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_io__storeAddrMisaligned; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_DTLBPF; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_DTLBENABLE; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_ISAMO2; // @[UnpipelinedLSU.scala 47:28]
  wire [63:0] lsExecUnit_io_in_bits_src1; // @[UnpipelinedLSU.scala 47:28]
  wire  lsExecUnit_DTLBFINISH; // @[UnpipelinedLSU.scala 47:28]
  wire [63:0] atomALU_io_src1; // @[UnpipelinedLSU.scala 98:25]
  wire [63:0] atomALU_io_src2; // @[UnpipelinedLSU.scala 98:25]
  wire [6:0] atomALU_io_func; // @[UnpipelinedLSU.scala 98:25]
  wire  atomALU_io_isWordOp; // @[UnpipelinedLSU.scala 98:25]
  wire [63:0] atomALU_io_result; // @[UnpipelinedLSU.scala 98:25]
  wire  atomReq = io__in_valid & io__in_bits_func[5]; // @[UnpipelinedLSU.scala 53:26]
  wire  _T_8 = io__in_bits_func == 7'h20; // @[LSU.scala 57:37]
  wire  _T_9 = ~_T_8; // @[LSU.scala 59:49]
  wire  _T_10 = io__in_bits_func[5] & _T_9; // @[LSU.scala 59:46]
  wire  _T_11 = io__in_bits_func == 7'h21; // @[LSU.scala 58:37]
  wire  _T_12 = ~_T_11; // @[LSU.scala 59:64]
  wire  _T_13 = _T_10 & _T_12; // @[LSU.scala 59:61]
  wire  amoReq = io__in_valid & _T_13; // @[UnpipelinedLSU.scala 54:26]
  wire  lrReq = io__in_valid & _T_8; // @[UnpipelinedLSU.scala 55:25]
  wire  scReq = io__in_valid & _T_11; // @[UnpipelinedLSU.scala 56:25]
  wire [2:0] funct3 = io__instr[14:12]; // @[UnpipelinedLSU.scala 64:26]
  wire  _T_17 = io__in_bits_src1 == lr_addr; // @[UnpipelinedLSU.scala 81:28]
  wire  _T_18 = ~_T_17; // @[UnpipelinedLSU.scala 81:21]
  wire  scInvalid = _T_18 & scReq; // @[UnpipelinedLSU.scala 81:40]
  reg [2:0] state; // @[UnpipelinedLSU.scala 95:24]
  reg [63:0] atomMemReg; // @[UnpipelinedLSU.scala 96:25]
  reg [63:0] atomRegReg; // @[UnpipelinedLSU.scala 97:25]
  wire  _T_19 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_22 = ~atomReq; // @[UnpipelinedLSU.scala 141:56]
  wire  _T_23 = io__in_valid & _T_22; // @[UnpipelinedLSU.scala 141:53]
  wire [63:0] _T_25 = io__in_bits_src1 + io__in_bits_src2; // @[UnpipelinedLSU.scala 143:46]
  wire  _T_26 = lsExecUnit_io__out_ready & lsExecUnit_io__out_valid; // @[Decoupled.scala 40:37]
  wire  _T_28 = lsExecUnit_io__out_valid | scInvalid; // @[UnpipelinedLSU.scala 148:66]
  wire  _T_30 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_33 = ~amoReq; // @[UnpipelinedLSU.scala 167:28]
  wire  _T_34 = _T_22 | _T_33; // @[UnpipelinedLSU.scala 167:25]
  wire  _T_35 = ~lrReq; // @[UnpipelinedLSU.scala 167:39]
  wire  _T_36 = _T_34 | _T_35; // @[UnpipelinedLSU.scala 167:36]
  wire  _T_37 = ~scReq; // @[UnpipelinedLSU.scala 167:49]
  wire  _T_38 = _T_36 | _T_37; // @[UnpipelinedLSU.scala 167:46]
  wire  _T_40 = _T_38 | reset; // @[UnpipelinedLSU.scala 167:15]
  wire  _T_41 = ~_T_40; // @[UnpipelinedLSU.scala 167:15]
  wire  _T_43 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire [1:0] _T_44 = funct3[0] ? 2'h3 : 2'h2; // @[UnpipelinedLSU.scala 188:42]
  wire  _T_55 = 3'h6 == state; // @[Conditional.scala 37:30]
  wire  _T_65 = 3'h7 == state; // @[Conditional.scala 37:30]
  wire [3:0] _T_66 = funct3[0] ? 4'hb : 4'ha; // @[UnpipelinedLSU.scala 219:42]
  wire  _T_79 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_93 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire [63:0] _GEN_11 = io__in_bits_src1; // @[Conditional.scala 39:67]
  wire  _GEN_14 = _T_93 & _T_26; // @[Conditional.scala 39:67]
  wire  _GEN_17 = _T_79 | _T_93; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_20 = _T_79 ? {{2'd0}, _T_44} : _T_66; // @[Conditional.scala 39:67]
  wire  _GEN_22 = _T_79 ? _T_26 : _GEN_14; // @[Conditional.scala 39:67]
  wire  _GEN_25 = _T_65 | _GEN_17; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_28 = _T_65 ? _T_66 : _GEN_20; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_29 = _T_65 ? atomMemReg : io__wdata; // @[Conditional.scala 39:67]
  wire  _GEN_30 = _T_65 ? _T_26 : _GEN_22; // @[Conditional.scala 39:67]
  wire  _GEN_33 = _T_55 ? 1'h0 : _GEN_25; // @[Conditional.scala 39:67]
  wire  _GEN_34 = _T_55 ? 1'h0 : 1'h1; // @[Conditional.scala 39:67]
  wire  _GEN_38 = _T_55 ? 1'h0 : _GEN_30; // @[Conditional.scala 39:67]
  wire  _GEN_42 = _T_43 | _GEN_33; // @[Conditional.scala 39:67]
  wire  _GEN_43 = _T_43 | _GEN_34; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_45 = _T_43 ? {{2'd0}, _T_44} : _GEN_28; // @[Conditional.scala 39:67]
  wire  _GEN_47 = _T_43 ? 1'h0 : _GEN_38; // @[Conditional.scala 39:67]
  wire  _GEN_52 = _T_30 | _GEN_42; // @[Conditional.scala 39:67]
  wire  _GEN_53 = _T_30 | _GEN_43; // @[Conditional.scala 39:67]
  wire [6:0] _GEN_55 = _T_30 ? io__in_bits_func : {{3'd0}, _GEN_45}; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_56 = _T_30 ? io__wdata : _GEN_29; // @[Conditional.scala 39:67]
  wire  _GEN_58 = _T_30 ? lsExecUnit_io__out_valid : _GEN_47; // @[Conditional.scala 39:67]
  wire  _GEN_68 = _T_19 ? _T_28 : _GEN_58; // @[Conditional.scala 40:58]
  wire  _T_107 = DTLBPF | io__loadAddrMisaligned; // @[UnpipelinedLSU.scala 257:17]
  wire  _T_108 = _T_107 | io__storeAddrMisaligned; // @[UnpipelinedLSU.scala 257:42]
  wire  _T_120 = lrReq | scReq; // @[UnpipelinedLSU.scala 270:38]
  wire  _T_121 = io__out_valid & _T_120; // @[UnpipelinedLSU.scala 270:28]
  wire  _T_122 = state == 3'h7; // @[UnpipelinedLSU.scala 275:52]
  wire [63:0] _T_123 = _T_122 ? atomRegReg : lsExecUnit_io__out_bits; // @[UnpipelinedLSU.scala 275:45]
  wire  setLr = _T_121; // @[UnpipelinedLSU.scala 70:21 UnpipelinedLSU.scala 270:11]
  wire  setLrVal = lrReq; // @[UnpipelinedLSU.scala 71:24 UnpipelinedLSU.scala 271:14]
  wire [63:0] setLrAddr = io__in_bits_src1; // @[UnpipelinedLSU.scala 72:25 UnpipelinedLSU.scala 272:15]
  wire  _GEN_77 = ~_T_19; // @[UnpipelinedLSU.scala 167:15]
  wire  _GEN_78 = _GEN_77 & _T_30; // @[UnpipelinedLSU.scala 167:15]
  LSExecUnit lsExecUnit ( // @[UnpipelinedLSU.scala 47:28]
    .clock(lsExecUnit_clock),
    .reset(lsExecUnit_reset),
    .io__in_valid(lsExecUnit_io__in_valid),
    .io__in_bits_src1(lsExecUnit_io__in_bits_src1),
    .io__in_bits_func(lsExecUnit_io__in_bits_func),
    .io__out_ready(lsExecUnit_io__out_ready),
    .io__out_valid(lsExecUnit_io__out_valid),
    .io__out_bits(lsExecUnit_io__out_bits),
    .io__wdata(lsExecUnit_io__wdata),
    .io__dmem_req_ready(lsExecUnit_io__dmem_req_ready),
    .io__dmem_req_valid(lsExecUnit_io__dmem_req_valid),
    .io__dmem_req_bits_addr(lsExecUnit_io__dmem_req_bits_addr),
    .io__dmem_req_bits_size(lsExecUnit_io__dmem_req_bits_size),
    .io__dmem_req_bits_cmd(lsExecUnit_io__dmem_req_bits_cmd),
    .io__dmem_req_bits_wmask(lsExecUnit_io__dmem_req_bits_wmask),
    .io__dmem_req_bits_wdata(lsExecUnit_io__dmem_req_bits_wdata),
    .io__dmem_resp_ready(lsExecUnit_io__dmem_resp_ready),
    .io__dmem_resp_valid(lsExecUnit_io__dmem_resp_valid),
    .io__dmem_resp_bits_rdata(lsExecUnit_io__dmem_resp_bits_rdata),
    .io__isMMIO(lsExecUnit_io__isMMIO),
    .io__dtlbPF(lsExecUnit_io__dtlbPF),
    .io__loadAddrMisaligned(lsExecUnit_io__loadAddrMisaligned),
    .io__storeAddrMisaligned(lsExecUnit_io__storeAddrMisaligned),
    .DTLBPF(lsExecUnit_DTLBPF),
    .DTLBENABLE(lsExecUnit_DTLBENABLE),
    .ISAMO2(lsExecUnit_ISAMO2),
    .io_in_bits_src1(lsExecUnit_io_in_bits_src1),
    .DTLBFINISH(lsExecUnit_DTLBFINISH)
  );
  AtomALU atomALU ( // @[UnpipelinedLSU.scala 98:25]
    .io_src1(atomALU_io_src1),
    .io_src2(atomALU_io_src2),
    .io_func(atomALU_io_func),
    .io_isWordOp(atomALU_io_isWordOp),
    .io_result(atomALU_io_result)
  );
  assign io__out_valid = _T_108 | _GEN_68; // @[UnpipelinedLSU.scala 125:32 UnpipelinedLSU.scala 137:36 UnpipelinedLSU.scala 148:38 UnpipelinedLSU.scala 166:36 UnpipelinedLSU.scala 191:36 UnpipelinedLSU.scala 208:36 UnpipelinedLSU.scala 222:36 UnpipelinedLSU.scala 236:36 UnpipelinedLSU.scala 250:36 UnpipelinedLSU.scala 259:20]
  assign io__out_bits = scReq ? {{63'd0}, scInvalid} : _T_123; // @[UnpipelinedLSU.scala 275:17]
  assign io__dmem_req_valid = lsExecUnit_io__dmem_req_valid; // @[UnpipelinedLSU.scala 274:13]
  assign io__dmem_req_bits_addr = lsExecUnit_io__dmem_req_bits_addr; // @[UnpipelinedLSU.scala 274:13]
  assign io__dmem_req_bits_size = lsExecUnit_io__dmem_req_bits_size; // @[UnpipelinedLSU.scala 274:13]
  assign io__dmem_req_bits_cmd = lsExecUnit_io__dmem_req_bits_cmd; // @[UnpipelinedLSU.scala 274:13]
  assign io__dmem_req_bits_wmask = lsExecUnit_io__dmem_req_bits_wmask; // @[UnpipelinedLSU.scala 274:13]
  assign io__dmem_req_bits_wdata = lsExecUnit_io__dmem_req_bits_wdata; // @[UnpipelinedLSU.scala 274:13]
  assign io__dtlbPF = lsExecUnit_io__dtlbPF; // @[UnpipelinedLSU.scala 49:15]
  assign io__loadAddrMisaligned = lsExecUnit_io__loadAddrMisaligned; // @[UnpipelinedLSU.scala 285:27]
  assign io__storeAddrMisaligned = lsExecUnit_io__storeAddrMisaligned; // @[UnpipelinedLSU.scala 286:28]
  assign setLr_0 = setLr;
  assign amoReq_0 = amoReq;
  assign io_in_bits_src1 = lsExecUnit_io_in_bits_src1;
  assign setLrAddr_0 = _GEN_11;
  assign setLrVal_0 = setLrVal;
  assign lsExecUnit_clock = clock;
  assign lsExecUnit_reset = reset;
  assign lsExecUnit_io__in_valid = _T_19 ? _T_23 : _GEN_52; // @[UnpipelinedLSU.scala 119:32 UnpipelinedLSU.scala 130:36 UnpipelinedLSU.scala 141:38 UnpipelinedLSU.scala 159:36 UnpipelinedLSU.scala 184:36 UnpipelinedLSU.scala 201:36 UnpipelinedLSU.scala 215:36 UnpipelinedLSU.scala 229:36 UnpipelinedLSU.scala 243:36]
  assign lsExecUnit_io__in_bits_src1 = _T_19 ? _T_25 : io__in_bits_src1; // @[UnpipelinedLSU.scala 143:38 UnpipelinedLSU.scala 186:36 UnpipelinedLSU.scala 217:36 UnpipelinedLSU.scala 231:36 UnpipelinedLSU.scala 245:36]
  assign lsExecUnit_io__in_bits_func = _T_19 ? io__in_bits_func : _GEN_55; // @[UnpipelinedLSU.scala 145:38 UnpipelinedLSU.scala 163:36 UnpipelinedLSU.scala 188:36 UnpipelinedLSU.scala 219:36 UnpipelinedLSU.scala 233:36 UnpipelinedLSU.scala 247:36]
  assign lsExecUnit_io__out_ready = _T_19 | _GEN_53; // @[UnpipelinedLSU.scala 142:38 UnpipelinedLSU.scala 160:36 UnpipelinedLSU.scala 185:36 UnpipelinedLSU.scala 202:36 UnpipelinedLSU.scala 216:36 UnpipelinedLSU.scala 230:36 UnpipelinedLSU.scala 244:36]
  assign lsExecUnit_io__wdata = _T_19 ? io__wdata : _GEN_56; // @[UnpipelinedLSU.scala 146:38 UnpipelinedLSU.scala 164:36 UnpipelinedLSU.scala 220:36 UnpipelinedLSU.scala 248:36]
  assign lsExecUnit_io__dmem_req_ready = io__dmem_req_ready; // @[UnpipelinedLSU.scala 274:13]
  assign lsExecUnit_io__dmem_resp_valid = io__dmem_resp_valid; // @[UnpipelinedLSU.scala 274:13]
  assign lsExecUnit_io__dmem_resp_bits_rdata = io__dmem_resp_bits_rdata; // @[UnpipelinedLSU.scala 274:13]
  assign lsExecUnit_DTLBPF = DTLBPF;
  assign lsExecUnit_DTLBENABLE = DTLBENABLE;
  assign lsExecUnit_ISAMO2 = amoReq;
  assign lsExecUnit_DTLBFINISH = DTLBFINISH;
  assign atomALU_io_src1 = atomMemReg; // @[UnpipelinedLSU.scala 99:21]
  assign atomALU_io_src2 = io__wdata; // @[UnpipelinedLSU.scala 100:21]
  assign atomALU_io_func = io__in_bits_func; // @[UnpipelinedLSU.scala 101:21]
  assign atomALU_io_isWordOp = ~funct3[0]; // @[UnpipelinedLSU.scala 102:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {2{`RANDOM}};
  atomMemReg = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  atomRegReg = _RAND_2[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 3'h0;
    end else if (_T_108) begin
      state <= 3'h0;
    end else if (_T_19) begin
      if (scReq) begin
        if (scInvalid) begin
          state <= 3'h0;
        end else begin
          state <= 3'h4;
        end
      end else if (lrReq) begin
        state <= 3'h3;
      end else if (amoReq) begin
        state <= 3'h5;
      end else begin
        state <= 3'h0;
      end
    end else if (_T_30) begin
      if (io__out_valid) begin
        state <= 3'h0;
      end
    end else if (_T_43) begin
      if (_T_26) begin
        state <= 3'h6;
      end
    end else if (_T_55) begin
      state <= 3'h7;
    end else if (_T_65) begin
      if (_T_26) begin
        state <= 3'h0;
      end
    end else if (_T_79) begin
      if (_T_26) begin
        state <= 3'h0;
      end
    end else if (_T_93) begin
      if (_T_26) begin
        state <= 3'h0;
      end
    end
    if (!(_T_19)) begin
      if (!(_T_30)) begin
        if (_T_43) begin
          atomMemReg <= lsExecUnit_io__out_bits;
        end else if (_T_55) begin
          atomMemReg <= atomALU_io_result;
        end
      end
    end
    if (!(_T_19)) begin
      if (!(_T_30)) begin
        if (_T_43) begin
          atomRegReg <= lsExecUnit_io__out_bits;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_GEN_78 & _T_41) begin
          $fwrite(32'h80000002,"Assertion failed\n    at UnpipelinedLSU.scala:167 assert(!atomReq || !amoReq || !lrReq || !scReq)\n"); // @[UnpipelinedLSU.scala 167:15]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_GEN_78 & _T_41) begin
          $fatal; // @[UnpipelinedLSU.scala 167:15]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Multiplier(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [64:0]  io_in_bits_0,
  input  [64:0]  io_in_bits_1,
  input          io_out_ready,
  output         io_out_valid,
  output [129:0] io_out_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [95:0] _RAND_0;
  reg [95:0] _RAND_1;
  reg [159:0] _RAND_2;
  reg [159:0] _RAND_3;
  reg [159:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  reg [64:0] _T; // @[MDU.scala 56:43]
  reg [64:0] _T_2; // @[MDU.scala 56:43]
  reg [129:0] _T_4; // @[MDU.scala 57:60]
  reg [129:0] _T_5; // @[MDU.scala 57:52]
  reg [129:0] _T_6; // @[MDU.scala 57:44]
  reg  _T_9; // @[MDU.scala 56:43]
  reg  _T_10; // @[MDU.scala 57:60]
  reg  _T_11; // @[MDU.scala 57:52]
  reg  _T_12; // @[MDU.scala 57:44]
  reg  busy; // @[MDU.scala 62:21]
  wire  _T_13 = ~busy; // @[MDU.scala 63:24]
  wire  _T_14 = io_in_valid & _T_13; // @[MDU.scala 63:21]
  wire  _GEN_0 = _T_14 | busy; // @[MDU.scala 63:31]
  assign io_in_ready = ~busy; // @[MDU.scala 65:15]
  assign io_out_valid = _T_12; // @[MDU.scala 60:16]
  assign io_out_bits = _T_6; // @[MDU.scala 59:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {3{`RANDOM}};
  _T = _RAND_0[64:0];
  _RAND_1 = {3{`RANDOM}};
  _T_2 = _RAND_1[64:0];
  _RAND_2 = {5{`RANDOM}};
  _T_4 = _RAND_2[129:0];
  _RAND_3 = {5{`RANDOM}};
  _T_5 = _RAND_3[129:0];
  _RAND_4 = {5{`RANDOM}};
  _T_6 = _RAND_4[129:0];
  _RAND_5 = {1{`RANDOM}};
  _T_9 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_10 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_11 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_12 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  busy = _RAND_9[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T <= io_in_bits_0;
    _T_2 <= io_in_bits_1;
    _T_4 <= $signed(_T) * $signed(_T_2);
    _T_5 <= _T_4;
    _T_6 <= _T_5;
    _T_9 <= io_in_ready & io_in_valid;
    _T_10 <= _T_9;
    _T_11 <= _T_10;
    _T_12 <= _T_11;
    if (reset) begin
      busy <= 1'h0;
    end else if (io_out_valid) begin
      busy <= 1'h0;
    end else begin
      busy <= _GEN_0;
    end
  end
endmodule
module Divider(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [63:0]  io_in_bits_0,
  input  [63:0]  io_in_bits_1,
  input          io_sign,
  output         io_out_valid,
  output [127:0] io_out_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [159:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [95:0] _RAND_5;
  reg [31:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[MDU.scala 77:22]
  wire  _T = state == 3'h0; // @[MDU.scala 78:23]
  wire  _T_1 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire  newReq = _T & _T_1; // @[MDU.scala 78:35]
  wire  divBy0 = io_in_bits_1 == 64'h0; // @[MDU.scala 81:18]
  reg [128:0] shiftReg; // @[MDU.scala 83:21]
  wire [64:0] hi = shiftReg[128:64]; // @[MDU.scala 84:20]
  wire [63:0] lo = shiftReg[63:0]; // @[MDU.scala 85:20]
  wire  aSign = io_in_bits_0[63] & io_sign; // @[MDU.scala 72:24]
  wire [63:0] _T_4 = 64'h0 - io_in_bits_0; // @[MDU.scala 73:16]
  wire [63:0] aVal = aSign ? _T_4 : io_in_bits_0; // @[MDU.scala 73:12]
  wire  bSign = io_in_bits_1[63] & io_sign; // @[MDU.scala 72:24]
  wire [63:0] _T_7 = 64'h0 - io_in_bits_1; // @[MDU.scala 73:16]
  reg  aSignReg; // @[Reg.scala 15:16]
  wire  _T_8 = aSign ^ bSign; // @[MDU.scala 90:35]
  wire  _T_9 = ~divBy0; // @[MDU.scala 90:47]
  wire  _T_10 = _T_8 & _T_9; // @[MDU.scala 90:44]
  reg  qSignReg; // @[Reg.scala 15:16]
  reg [63:0] bReg; // @[Reg.scala 15:16]
  wire [64:0] _T_11 = {aVal,1'h0}; // @[Cat.scala 29:58]
  reg [64:0] aValx2Reg; // @[Reg.scala 15:16]
  reg [5:0] value; // @[Counter.scala 29:33]
  wire  _T_12 = state == 3'h1; // @[MDU.scala 97:22]
  wire  _T_15 = |bReg[63:32]; // @[CircuitMath.scala 37:22]
  wire  _T_18 = |bReg[63:48]; // @[CircuitMath.scala 37:22]
  wire  _T_21 = |bReg[63:56]; // @[CircuitMath.scala 37:22]
  wire  _T_24 = |bReg[63:60]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_28 = bReg[62] ? 2'h2 : {{1'd0}, bReg[61]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_29 = bReg[63] ? 2'h3 : _T_28; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_33 = bReg[58] ? 2'h2 : {{1'd0}, bReg[57]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_34 = bReg[59] ? 2'h3 : _T_33; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_35 = _T_24 ? _T_29 : _T_34; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_36 = {_T_24,_T_35}; // @[Cat.scala 29:58]
  wire  _T_39 = |bReg[55:52]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_43 = bReg[54] ? 2'h2 : {{1'd0}, bReg[53]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_44 = bReg[55] ? 2'h3 : _T_43; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_48 = bReg[50] ? 2'h2 : {{1'd0}, bReg[49]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_49 = bReg[51] ? 2'h3 : _T_48; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_50 = _T_39 ? _T_44 : _T_49; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_51 = {_T_39,_T_50}; // @[Cat.scala 29:58]
  wire [2:0] _T_52 = _T_21 ? _T_36 : _T_51; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_53 = {_T_21,_T_52}; // @[Cat.scala 29:58]
  wire  _T_56 = |bReg[47:40]; // @[CircuitMath.scala 37:22]
  wire  _T_59 = |bReg[47:44]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_63 = bReg[46] ? 2'h2 : {{1'd0}, bReg[45]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_64 = bReg[47] ? 2'h3 : _T_63; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_68 = bReg[42] ? 2'h2 : {{1'd0}, bReg[41]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_69 = bReg[43] ? 2'h3 : _T_68; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_70 = _T_59 ? _T_64 : _T_69; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_71 = {_T_59,_T_70}; // @[Cat.scala 29:58]
  wire  _T_74 = |bReg[39:36]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_78 = bReg[38] ? 2'h2 : {{1'd0}, bReg[37]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_79 = bReg[39] ? 2'h3 : _T_78; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_83 = bReg[34] ? 2'h2 : {{1'd0}, bReg[33]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_84 = bReg[35] ? 2'h3 : _T_83; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_85 = _T_74 ? _T_79 : _T_84; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_86 = {_T_74,_T_85}; // @[Cat.scala 29:58]
  wire [2:0] _T_87 = _T_56 ? _T_71 : _T_86; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_88 = {_T_56,_T_87}; // @[Cat.scala 29:58]
  wire [3:0] _T_89 = _T_18 ? _T_53 : _T_88; // @[CircuitMath.scala 38:21]
  wire [4:0] _T_90 = {_T_18,_T_89}; // @[Cat.scala 29:58]
  wire  _T_93 = |bReg[31:16]; // @[CircuitMath.scala 37:22]
  wire  _T_96 = |bReg[31:24]; // @[CircuitMath.scala 37:22]
  wire  _T_99 = |bReg[31:28]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_103 = bReg[30] ? 2'h2 : {{1'd0}, bReg[29]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_104 = bReg[31] ? 2'h3 : _T_103; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_108 = bReg[26] ? 2'h2 : {{1'd0}, bReg[25]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_109 = bReg[27] ? 2'h3 : _T_108; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_110 = _T_99 ? _T_104 : _T_109; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_111 = {_T_99,_T_110}; // @[Cat.scala 29:58]
  wire  _T_114 = |bReg[23:20]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_118 = bReg[22] ? 2'h2 : {{1'd0}, bReg[21]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_119 = bReg[23] ? 2'h3 : _T_118; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_123 = bReg[18] ? 2'h2 : {{1'd0}, bReg[17]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_124 = bReg[19] ? 2'h3 : _T_123; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_125 = _T_114 ? _T_119 : _T_124; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_126 = {_T_114,_T_125}; // @[Cat.scala 29:58]
  wire [2:0] _T_127 = _T_96 ? _T_111 : _T_126; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_128 = {_T_96,_T_127}; // @[Cat.scala 29:58]
  wire  _T_131 = |bReg[15:8]; // @[CircuitMath.scala 37:22]
  wire  _T_134 = |bReg[15:12]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_138 = bReg[14] ? 2'h2 : {{1'd0}, bReg[13]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_139 = bReg[15] ? 2'h3 : _T_138; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_143 = bReg[10] ? 2'h2 : {{1'd0}, bReg[9]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_144 = bReg[11] ? 2'h3 : _T_143; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_145 = _T_134 ? _T_139 : _T_144; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_146 = {_T_134,_T_145}; // @[Cat.scala 29:58]
  wire  _T_149 = |bReg[7:4]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_153 = bReg[6] ? 2'h2 : {{1'd0}, bReg[5]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_154 = bReg[7] ? 2'h3 : _T_153; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_158 = bReg[2] ? 2'h2 : {{1'd0}, bReg[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_159 = bReg[3] ? 2'h3 : _T_158; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_160 = _T_149 ? _T_154 : _T_159; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_161 = {_T_149,_T_160}; // @[Cat.scala 29:58]
  wire [2:0] _T_162 = _T_131 ? _T_146 : _T_161; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_163 = {_T_131,_T_162}; // @[Cat.scala 29:58]
  wire [3:0] _T_164 = _T_93 ? _T_128 : _T_163; // @[CircuitMath.scala 38:21]
  wire [4:0] _T_165 = {_T_93,_T_164}; // @[Cat.scala 29:58]
  wire [4:0] _T_166 = _T_15 ? _T_90 : _T_165; // @[CircuitMath.scala 38:21]
  wire [5:0] _T_167 = {_T_15,_T_166}; // @[Cat.scala 29:58]
  wire [6:0] _GEN_18 = {{1'd0}, _T_167}; // @[MDU.scala 105:31]
  wire [6:0] _T_168 = 7'h40 | _GEN_18; // @[MDU.scala 105:31]
  wire  _T_171 = |aValx2Reg[64]; // @[CircuitMath.scala 37:22]
  wire  _T_174 = |aValx2Reg[63:32]; // @[CircuitMath.scala 37:22]
  wire  _T_177 = |aValx2Reg[63:48]; // @[CircuitMath.scala 37:22]
  wire  _T_180 = |aValx2Reg[63:56]; // @[CircuitMath.scala 37:22]
  wire  _T_183 = |aValx2Reg[63:60]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_187 = aValx2Reg[62] ? 2'h2 : {{1'd0}, aValx2Reg[61]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_188 = aValx2Reg[63] ? 2'h3 : _T_187; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_192 = aValx2Reg[58] ? 2'h2 : {{1'd0}, aValx2Reg[57]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_193 = aValx2Reg[59] ? 2'h3 : _T_192; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_194 = _T_183 ? _T_188 : _T_193; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_195 = {_T_183,_T_194}; // @[Cat.scala 29:58]
  wire  _T_198 = |aValx2Reg[55:52]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_202 = aValx2Reg[54] ? 2'h2 : {{1'd0}, aValx2Reg[53]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_203 = aValx2Reg[55] ? 2'h3 : _T_202; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_207 = aValx2Reg[50] ? 2'h2 : {{1'd0}, aValx2Reg[49]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_208 = aValx2Reg[51] ? 2'h3 : _T_207; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_209 = _T_198 ? _T_203 : _T_208; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_210 = {_T_198,_T_209}; // @[Cat.scala 29:58]
  wire [2:0] _T_211 = _T_180 ? _T_195 : _T_210; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_212 = {_T_180,_T_211}; // @[Cat.scala 29:58]
  wire  _T_215 = |aValx2Reg[47:40]; // @[CircuitMath.scala 37:22]
  wire  _T_218 = |aValx2Reg[47:44]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_222 = aValx2Reg[46] ? 2'h2 : {{1'd0}, aValx2Reg[45]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_223 = aValx2Reg[47] ? 2'h3 : _T_222; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_227 = aValx2Reg[42] ? 2'h2 : {{1'd0}, aValx2Reg[41]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_228 = aValx2Reg[43] ? 2'h3 : _T_227; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_229 = _T_218 ? _T_223 : _T_228; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_230 = {_T_218,_T_229}; // @[Cat.scala 29:58]
  wire  _T_233 = |aValx2Reg[39:36]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_237 = aValx2Reg[38] ? 2'h2 : {{1'd0}, aValx2Reg[37]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_238 = aValx2Reg[39] ? 2'h3 : _T_237; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_242 = aValx2Reg[34] ? 2'h2 : {{1'd0}, aValx2Reg[33]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_243 = aValx2Reg[35] ? 2'h3 : _T_242; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_244 = _T_233 ? _T_238 : _T_243; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_245 = {_T_233,_T_244}; // @[Cat.scala 29:58]
  wire [2:0] _T_246 = _T_215 ? _T_230 : _T_245; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_247 = {_T_215,_T_246}; // @[Cat.scala 29:58]
  wire [3:0] _T_248 = _T_177 ? _T_212 : _T_247; // @[CircuitMath.scala 38:21]
  wire [4:0] _T_249 = {_T_177,_T_248}; // @[Cat.scala 29:58]
  wire  _T_252 = |aValx2Reg[31:16]; // @[CircuitMath.scala 37:22]
  wire  _T_255 = |aValx2Reg[31:24]; // @[CircuitMath.scala 37:22]
  wire  _T_258 = |aValx2Reg[31:28]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_262 = aValx2Reg[30] ? 2'h2 : {{1'd0}, aValx2Reg[29]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_263 = aValx2Reg[31] ? 2'h3 : _T_262; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_267 = aValx2Reg[26] ? 2'h2 : {{1'd0}, aValx2Reg[25]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_268 = aValx2Reg[27] ? 2'h3 : _T_267; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_269 = _T_258 ? _T_263 : _T_268; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_270 = {_T_258,_T_269}; // @[Cat.scala 29:58]
  wire  _T_273 = |aValx2Reg[23:20]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_277 = aValx2Reg[22] ? 2'h2 : {{1'd0}, aValx2Reg[21]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_278 = aValx2Reg[23] ? 2'h3 : _T_277; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_282 = aValx2Reg[18] ? 2'h2 : {{1'd0}, aValx2Reg[17]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_283 = aValx2Reg[19] ? 2'h3 : _T_282; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_284 = _T_273 ? _T_278 : _T_283; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_285 = {_T_273,_T_284}; // @[Cat.scala 29:58]
  wire [2:0] _T_286 = _T_255 ? _T_270 : _T_285; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_287 = {_T_255,_T_286}; // @[Cat.scala 29:58]
  wire  _T_290 = |aValx2Reg[15:8]; // @[CircuitMath.scala 37:22]
  wire  _T_293 = |aValx2Reg[15:12]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_297 = aValx2Reg[14] ? 2'h2 : {{1'd0}, aValx2Reg[13]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_298 = aValx2Reg[15] ? 2'h3 : _T_297; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_302 = aValx2Reg[10] ? 2'h2 : {{1'd0}, aValx2Reg[9]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_303 = aValx2Reg[11] ? 2'h3 : _T_302; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_304 = _T_293 ? _T_298 : _T_303; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_305 = {_T_293,_T_304}; // @[Cat.scala 29:58]
  wire  _T_308 = |aValx2Reg[7:4]; // @[CircuitMath.scala 37:22]
  wire [1:0] _T_312 = aValx2Reg[6] ? 2'h2 : {{1'd0}, aValx2Reg[5]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_313 = aValx2Reg[7] ? 2'h3 : _T_312; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_317 = aValx2Reg[2] ? 2'h2 : {{1'd0}, aValx2Reg[1]}; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_318 = aValx2Reg[3] ? 2'h3 : _T_317; // @[CircuitMath.scala 32:10]
  wire [1:0] _T_319 = _T_308 ? _T_313 : _T_318; // @[CircuitMath.scala 38:21]
  wire [2:0] _T_320 = {_T_308,_T_319}; // @[Cat.scala 29:58]
  wire [2:0] _T_321 = _T_290 ? _T_305 : _T_320; // @[CircuitMath.scala 38:21]
  wire [3:0] _T_322 = {_T_290,_T_321}; // @[Cat.scala 29:58]
  wire [3:0] _T_323 = _T_252 ? _T_287 : _T_322; // @[CircuitMath.scala 38:21]
  wire [4:0] _T_324 = {_T_252,_T_323}; // @[Cat.scala 29:58]
  wire [4:0] _T_325 = _T_174 ? _T_249 : _T_324; // @[CircuitMath.scala 38:21]
  wire [5:0] _T_326 = {_T_174,_T_325}; // @[Cat.scala 29:58]
  wire [5:0] _T_327 = _T_171 ? 6'h0 : _T_326; // @[CircuitMath.scala 38:21]
  wire [6:0] _T_328 = {_T_171,_T_327}; // @[Cat.scala 29:58]
  wire [6:0] _T_330 = _T_168 - _T_328; // @[MDU.scala 105:45]
  wire  _T_331 = _T_330 >= 7'h3f; // @[MDU.scala 109:52]
  wire [6:0] _T_332 = _T_331 ? 7'h3f : _T_330; // @[MDU.scala 109:38]
  wire [6:0] _T_333 = divBy0 ? 7'h0 : _T_332; // @[MDU.scala 109:21]
  wire  _T_334 = state == 3'h2; // @[MDU.scala 111:22]
  wire [127:0] _GEN_19 = {{63'd0}, aValx2Reg}; // @[MDU.scala 112:27]
  wire [127:0] _T_335 = _GEN_19 << value; // @[MDU.scala 112:27]
  wire  _T_336 = state == 3'h3; // @[MDU.scala 114:22]
  wire [64:0] _GEN_20 = {{1'd0}, bReg}; // @[MDU.scala 115:28]
  wire  _T_337 = hi >= _GEN_20; // @[MDU.scala 115:28]
  wire [64:0] _T_339 = hi - _GEN_20; // @[MDU.scala 116:36]
  wire [64:0] _T_340 = _T_337 ? _T_339 : hi; // @[MDU.scala 116:24]
  wire [128:0] _T_343 = {_T_340[63:0],lo,_T_337}; // @[Cat.scala 29:58]
  wire  _T_344 = value == 6'h3f; // @[Counter.scala 38:24]
  wire [5:0] _T_346 = value + 6'h1; // @[Counter.scala 39:22]
  wire  _T_348 = state == 3'h4; // @[MDU.scala 119:22]
  wire [5:0] _GEN_7 = _T_336 ? _T_346 : value; // @[MDU.scala 114:37]
  wire [5:0] _GEN_11 = _T_334 ? value : _GEN_7; // @[MDU.scala 111:35]
  wire [6:0] _GEN_12 = _T_12 ? _T_333 : {{1'd0}, _GEN_11}; // @[MDU.scala 97:34]
  wire [6:0] _GEN_16 = newReq ? {{1'd0}, value} : _GEN_12; // @[MDU.scala 95:17]
  wire [63:0] r = hi[64:1]; // @[MDU.scala 123:13]
  wire [63:0] _T_350 = 64'h0 - lo; // @[MDU.scala 124:28]
  wire [63:0] resQ = qSignReg ? _T_350 : lo; // @[MDU.scala 124:17]
  wire [63:0] _T_352 = 64'h0 - r; // @[MDU.scala 125:28]
  wire [63:0] resR = aSignReg ? _T_352 : r; // @[MDU.scala 125:17]
  assign io_in_ready = state == 3'h0; // @[MDU.scala 129:15]
  assign io_out_valid = state == 3'h4; // @[MDU.scala 128:16]
  assign io_out_bits = {resR,resQ}; // @[MDU.scala 126:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {5{`RANDOM}};
  shiftReg = _RAND_1[128:0];
  _RAND_2 = {1{`RANDOM}};
  aSignReg = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  qSignReg = _RAND_3[0:0];
  _RAND_4 = {2{`RANDOM}};
  bReg = _RAND_4[63:0];
  _RAND_5 = {3{`RANDOM}};
  aValx2Reg = _RAND_5[64:0];
  _RAND_6 = {1{`RANDOM}};
  value = _RAND_6[5:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 3'h0;
    end else if (newReq) begin
      state <= 3'h1;
    end else if (_T_12) begin
      state <= 3'h2;
    end else if (_T_334) begin
      state <= 3'h3;
    end else if (_T_336) begin
      if (_T_344) begin
        state <= 3'h4;
      end
    end else if (_T_348) begin
      state <= 3'h0;
    end
    if (!(newReq)) begin
      if (!(_T_12)) begin
        if (_T_334) begin
          shiftReg <= {{1'd0}, _T_335};
        end else if (_T_336) begin
          shiftReg <= _T_343;
        end
      end
    end
    if (newReq) begin
      aSignReg <= aSign;
    end
    if (newReq) begin
      qSignReg <= _T_10;
    end
    if (newReq) begin
      if (bSign) begin
        bReg <= _T_7;
      end else begin
        bReg <= io_in_bits_1;
      end
    end
    if (newReq) begin
      aValx2Reg <= _T_11;
    end
    if (reset) begin
      value <= 6'h0;
    end else begin
      value <= _GEN_16[5:0];
    end
  end
endmodule
module MDU(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [63:0] io_in_bits_src1,
  input  [63:0] io_in_bits_src2,
  input  [6:0]  io_in_bits_func,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
`endif // RANDOMIZE_REG_INIT
  wire  mul_clock; // @[MDU.scala 151:19]
  wire  mul_reset; // @[MDU.scala 151:19]
  wire  mul_io_in_ready; // @[MDU.scala 151:19]
  wire  mul_io_in_valid; // @[MDU.scala 151:19]
  wire [64:0] mul_io_in_bits_0; // @[MDU.scala 151:19]
  wire [64:0] mul_io_in_bits_1; // @[MDU.scala 151:19]
  wire  mul_io_out_ready; // @[MDU.scala 151:19]
  wire  mul_io_out_valid; // @[MDU.scala 151:19]
  wire [129:0] mul_io_out_bits; // @[MDU.scala 151:19]
  wire  div_clock; // @[MDU.scala 152:19]
  wire  div_reset; // @[MDU.scala 152:19]
  wire  div_io_in_ready; // @[MDU.scala 152:19]
  wire  div_io_in_valid; // @[MDU.scala 152:19]
  wire [63:0] div_io_in_bits_0; // @[MDU.scala 152:19]
  wire [63:0] div_io_in_bits_1; // @[MDU.scala 152:19]
  wire  div_io_sign; // @[MDU.scala 152:19]
  wire  div_io_out_valid; // @[MDU.scala 152:19]
  wire [127:0] div_io_out_bits; // @[MDU.scala 152:19]
  wire  isDiv = io_in_bits_func[2]; // @[MDU.scala 41:27]
  wire  _T_2 = ~io_in_bits_func[0]; // @[MDU.scala 42:42]
  wire  isDivSign = isDiv & _T_2; // @[MDU.scala 42:39]
  wire  isW = io_in_bits_func[3]; // @[MDU.scala 43:25]
  wire [64:0] _T_4 = {1'h0,io_in_bits_src1}; // @[Cat.scala 29:58]
  wire [64:0] _T_6 = {io_in_bits_src1[63],io_in_bits_src1}; // @[Cat.scala 29:58]
  wire  _T_10 = 2'h0 == io_in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_11 = 2'h1 == io_in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_12 = 2'h2 == io_in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire  _T_13 = 2'h3 == io_in_bits_func[1:0]; // @[LookupTree.scala 24:34]
  wire [64:0] _T_14 = _T_10 ? _T_4 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_15 = _T_11 ? _T_6 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_16 = _T_12 ? _T_6 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_17 = _T_13 ? _T_4 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_18 = _T_14 | _T_15; // @[Mux.scala 27:72]
  wire [64:0] _T_19 = _T_18 | _T_16; // @[Mux.scala 27:72]
  wire [64:0] _T_23 = {1'h0,io_in_bits_src2}; // @[Cat.scala 29:58]
  wire [64:0] _T_25 = {io_in_bits_src2[63],io_in_bits_src2}; // @[Cat.scala 29:58]
  wire [64:0] _T_32 = _T_10 ? _T_23 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_33 = _T_11 ? _T_25 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_34 = _T_12 ? _T_23 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_35 = _T_13 ? _T_23 : 65'h0; // @[Mux.scala 27:72]
  wire [64:0] _T_36 = _T_32 | _T_33; // @[Mux.scala 27:72]
  wire [64:0] _T_37 = _T_36 | _T_34; // @[Mux.scala 27:72]
  wire [31:0] _T_43 = io_in_bits_src1[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_44 = {_T_43,io_in_bits_src1[31:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_46 = {32'h0,io_in_bits_src1[31:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_47 = isDivSign ? _T_44 : _T_46; // @[MDU.scala 169:47]
  wire [31:0] _T_52 = io_in_bits_src2[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_53 = {_T_52,io_in_bits_src2[31:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_55 = {32'h0,io_in_bits_src2[31:0]}; // @[Cat.scala 29:58]
  wire [63:0] _T_56 = isDivSign ? _T_53 : _T_55; // @[MDU.scala 169:47]
  wire  _T_58 = ~isDiv; // @[MDU.scala 173:37]
  wire  _T_62 = io_in_bits_func[1:0] == 2'h0; // @[MDU.scala 176:30]
  wire [63:0] mulRes = _T_62 ? mul_io_out_bits[63:0] : mul_io_out_bits[127:64]; // @[MDU.scala 176:19]
  wire [63:0] divRes = io_in_bits_func[1] ? div_io_out_bits[127:64] : div_io_out_bits[63:0]; // @[MDU.scala 177:19]
  wire [63:0] res = isDiv ? divRes : mulRes; // @[MDU.scala 178:16]
  wire [31:0] _T_71 = res[31] ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_72 = {_T_71,res[31:0]}; // @[Cat.scala 29:58]
  wire  _T_74 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  reg  _T_75; // @[MDU.scala 181:50]
  wire  isDivReg = _T_74 ? isDiv : _T_75; // @[MDU.scala 181:21]
  wire  _T_87 = mul_io_out_ready & mul_io_out_valid; // @[Decoupled.scala 40:37]
  Multiplier mul ( // @[MDU.scala 151:19]
    .clock(mul_clock),
    .reset(mul_reset),
    .io_in_ready(mul_io_in_ready),
    .io_in_valid(mul_io_in_valid),
    .io_in_bits_0(mul_io_in_bits_0),
    .io_in_bits_1(mul_io_in_bits_1),
    .io_out_ready(mul_io_out_ready),
    .io_out_valid(mul_io_out_valid),
    .io_out_bits(mul_io_out_bits)
  );
  Divider div ( // @[MDU.scala 152:19]
    .clock(div_clock),
    .reset(div_reset),
    .io_in_ready(div_io_in_ready),
    .io_in_valid(div_io_in_valid),
    .io_in_bits_0(div_io_in_bits_0),
    .io_in_bits_1(div_io_in_bits_1),
    .io_sign(div_io_sign),
    .io_out_valid(div_io_out_valid),
    .io_out_bits(div_io_out_bits)
  );
  assign io_in_ready = isDiv ? div_io_in_ready : mul_io_in_ready; // @[MDU.scala 182:15]
  assign io_out_valid = isDivReg ? div_io_out_valid : mul_io_out_valid; // @[MDU.scala 183:16]
  assign io_out_bits = isW ? _T_72 : res; // @[MDU.scala 179:15]
  assign mul_clock = clock;
  assign mul_reset = reset;
  assign mul_io_in_valid = io_in_valid & _T_58; // @[MDU.scala 173:19]
  assign mul_io_in_bits_0 = _T_19 | _T_17; // @[MDU.scala 166:21]
  assign mul_io_in_bits_1 = _T_37 | _T_35; // @[MDU.scala 167:21]
  assign mul_io_out_ready = 1'h1; // @[MDU.scala 155:17]
  assign div_clock = clock;
  assign div_reset = reset;
  assign div_io_in_valid = io_in_valid & isDiv; // @[MDU.scala 174:19]
  assign div_io_in_bits_0 = isW ? _T_47 : io_in_bits_src1; // @[MDU.scala 170:21]
  assign div_io_in_bits_1 = isW ? _T_56 : io_in_bits_src2; // @[MDU.scala 171:21]
  assign div_io_sign = isDiv & _T_2; // @[MDU.scala 154:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_75 = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_75 <= io_in_bits_func[2];
  end
endmodule
module CSR(
  input         clock,
  input         reset,
  input         io_in_valid,
  input  [63:0] io_in_bits_src1,
  input  [63:0] io_in_bits_src2,
  input  [6:0]  io_in_bits_func,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits,
  input  [63:0] io_cfIn_instr,
  input  [38:0] io_cfIn_pc,
  input         io_cfIn_exceptionVec_1,
  input         io_cfIn_exceptionVec_2,
  input         io_cfIn_exceptionVec_4,
  input         io_cfIn_exceptionVec_6,
  input         io_cfIn_exceptionVec_12,
  input         io_cfIn_intrVec_0,
  input         io_cfIn_intrVec_1,
  input         io_cfIn_intrVec_2,
  input         io_cfIn_intrVec_3,
  input         io_cfIn_intrVec_4,
  input         io_cfIn_intrVec_5,
  input         io_cfIn_intrVec_6,
  input         io_cfIn_intrVec_7,
  input         io_cfIn_intrVec_8,
  input         io_cfIn_intrVec_9,
  input         io_cfIn_intrVec_10,
  input         io_cfIn_intrVec_11,
  input         io_cfIn_crossPageIPFFix,
  output [38:0] io_redirect_target,
  output        io_redirect_valid,
  input         io_instrValid,
  output [1:0]  io_imemMMU_priviledgeMode,
  output [1:0]  io_dmemMMU_priviledgeMode,
  output        io_dmemMMU_status_sum,
  output        io_dmemMMU_status_mxr,
  input         io_dmemMMU_loadPF,
  input         io_dmemMMU_storePF,
  input  [38:0] io_dmemMMU_addr,
  output        io_wenFix,
  input         set_lr,
  output [63:0] perfCnts_2_0,
  output [63:0] satp_0,
  input         perfCntCondMinstret,
  input         mtip_0,
  input         meip_0,
  input  [63:0] LSUADDR,
  output [11:0] intrVec_0,
  input         msip_0,
  input  [63:0] set_lr_addr,
  input         perfCntCondMultiCommit,
  input         set_lr_val,
  output [63:0] lrAddr_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [63:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [63:0] _RAND_12;
  reg [63:0] _RAND_13;
  reg [63:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [63:0] _RAND_16;
  reg [63:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [63:0] _RAND_32;
`endif // RANDOMIZE_REG_INIT
  reg [63:0] mtvec; // @[CSR.scala 251:22]
  reg [63:0] mcounteren; // @[CSR.scala 252:27]
  reg [63:0] mcause; // @[CSR.scala 253:23]
  reg [63:0] mtval; // @[CSR.scala 254:22]
  reg [63:0] mepc; // @[CSR.scala 255:17]
  reg [63:0] mie; // @[CSR.scala 257:20]
  reg [63:0] mipReg; // @[CSR.scala 259:24]
  wire [11:0] _T_23 = {meip_0,1'h0,1'h0,1'h0,mtip_0,1'h0,2'h0,msip_0,3'h0}; // @[CSR.scala 261:22]
  wire [63:0] _GEN_78 = {{52'd0}, _T_23}; // @[CSR.scala 261:29]
  wire [63:0] _T_24 = _GEN_78 | mipReg; // @[CSR.scala 261:29]
  wire  mip_s_u = _T_24[0]; // @[CSR.scala 261:47]
  wire  mip_s_s = _T_24[1]; // @[CSR.scala 261:47]
  wire  mip_s_h = _T_24[2]; // @[CSR.scala 261:47]
  wire  mip_s_m = _T_24[3]; // @[CSR.scala 261:47]
  wire  mip_t_u = _T_24[4]; // @[CSR.scala 261:47]
  wire  mip_t_s = _T_24[5]; // @[CSR.scala 261:47]
  wire  mip_t_h = _T_24[6]; // @[CSR.scala 261:47]
  wire  mip_t_m = _T_24[7]; // @[CSR.scala 261:47]
  wire  mip_e_u = _T_24[8]; // @[CSR.scala 261:47]
  wire  mip_e_s = _T_24[9]; // @[CSR.scala 261:47]
  wire  mip_e_h = _T_24[10]; // @[CSR.scala 261:47]
  wire  mip_e_m = _T_24[11]; // @[CSR.scala 261:47]
  reg [63:0] misa; // @[CSR.scala 269:21]
  reg [63:0] mstatus; // @[CSR.scala 277:24]
  wire  mstatusStruct_ie_u = mstatus[0]; // @[CSR.scala 298:39]
  wire  mstatusStruct_ie_s = mstatus[1]; // @[CSR.scala 298:39]
  wire  mstatusStruct_ie_h = mstatus[2]; // @[CSR.scala 298:39]
  wire  mstatusStruct_ie_m = mstatus[3]; // @[CSR.scala 298:39]
  wire  mstatusStruct_pie_u = mstatus[4]; // @[CSR.scala 298:39]
  wire  mstatusStruct_pie_s = mstatus[5]; // @[CSR.scala 298:39]
  wire  mstatusStruct_pie_h = mstatus[6]; // @[CSR.scala 298:39]
  wire  mstatusStruct_pie_m = mstatus[7]; // @[CSR.scala 298:39]
  wire  mstatusStruct_spp = mstatus[8]; // @[CSR.scala 298:39]
  wire [1:0] mstatusStruct_hpp = mstatus[10:9]; // @[CSR.scala 298:39]
  wire [1:0] mstatusStruct_mpp = mstatus[12:11]; // @[CSR.scala 298:39]
  wire [1:0] mstatusStruct_fs = mstatus[14:13]; // @[CSR.scala 298:39]
  wire [1:0] mstatusStruct_xs = mstatus[16:15]; // @[CSR.scala 298:39]
  wire  mstatusStruct_mprv = mstatus[17]; // @[CSR.scala 298:39]
  wire  mstatusStruct_sum = mstatus[18]; // @[CSR.scala 298:39]
  wire  mstatusStruct_mxr = mstatus[19]; // @[CSR.scala 298:39]
  wire  mstatusStruct_tvm = mstatus[20]; // @[CSR.scala 298:39]
  wire  mstatusStruct_tw = mstatus[21]; // @[CSR.scala 298:39]
  wire  mstatusStruct_tsr = mstatus[22]; // @[CSR.scala 298:39]
  wire [8:0] mstatusStruct_pad0 = mstatus[31:23]; // @[CSR.scala 298:39]
  wire [1:0] mstatusStruct_uxl = mstatus[33:32]; // @[CSR.scala 298:39]
  wire [1:0] mstatusStruct_sxl = mstatus[35:34]; // @[CSR.scala 298:39]
  wire [26:0] mstatusStruct_pad1 = mstatus[62:36]; // @[CSR.scala 298:39]
  wire  mstatusStruct_sd = mstatus[63]; // @[CSR.scala 298:39]
  reg [63:0] medeleg; // @[CSR.scala 305:24]
  reg [63:0] mideleg; // @[CSR.scala 306:24]
  reg [63:0] mscratch; // @[CSR.scala 307:25]
  reg [63:0] pmpcfg0; // @[CSR.scala 309:24]
  reg [63:0] pmpcfg1; // @[CSR.scala 310:24]
  reg [63:0] pmpcfg2; // @[CSR.scala 311:24]
  reg [63:0] pmpcfg3; // @[CSR.scala 312:24]
  reg [63:0] pmpaddr0; // @[CSR.scala 313:25]
  reg [63:0] pmpaddr1; // @[CSR.scala 314:25]
  reg [63:0] pmpaddr2; // @[CSR.scala 315:25]
  reg [63:0] pmpaddr3; // @[CSR.scala 316:25]
  reg [63:0] stvec; // @[CSR.scala 330:22]
  wire [63:0] sieMask = 64'h222 & mideleg; // @[CSR.scala 332:26]
  reg [63:0] satp; // @[CSR.scala 335:21]
  reg [63:0] sepc; // @[CSR.scala 336:21]
  reg [63:0] scause; // @[CSR.scala 337:23]
  reg [63:0] stval; // @[CSR.scala 338:18]
  reg [63:0] sscratch; // @[CSR.scala 339:25]
  reg [63:0] scounteren; // @[CSR.scala 340:27]
  reg  lr; // @[CSR.scala 353:19]
  reg [63:0] lrAddr; // @[CSR.scala 354:23]
  reg [1:0] priviledgeMode; // @[CSR.scala 367:31]
  reg [63:0] perfCnts_0; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_1; // @[CSR.scala 372:47]
  reg [63:0] perfCnts_2; // @[CSR.scala 372:47]
  wire [5:0] _T_107 = {mip_t_s,mip_t_u,mip_s_m,mip_s_h,mip_s_s,mip_s_u}; // @[CSR.scala 415:27]
  wire [11:0] _T_113 = {mip_e_m,mip_e_h,mip_e_s,mip_e_u,mip_t_m,mip_t_h,_T_107}; // @[CSR.scala 415:27]
  wire [11:0] addr = io_in_bits_src2[11:0]; // @[CSR.scala 455:18]
  wire [63:0] csri = {59'h0,io_cfIn_instr[19:15]}; // @[Cat.scala 29:58]
  wire  _T_257 = 12'hf12 == addr; // @[LookupTree.scala 24:34]
  wire  _T_258 = 12'h180 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_295 = _T_258 ? satp : 64'h0; // @[Mux.scala 27:72]
  wire  _T_259 = 12'h3b1 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_296 = _T_259 ? pmpaddr1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_332 = _T_295 | _T_296; // @[Mux.scala 27:72]
  wire  _T_260 = 12'h3a2 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_297 = _T_260 ? pmpcfg2 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_333 = _T_332 | _T_297; // @[Mux.scala 27:72]
  wire  _T_261 = 12'h140 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_298 = _T_261 ? sscratch : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_334 = _T_333 | _T_298; // @[Mux.scala 27:72]
  wire  _T_262 = 12'h302 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_299 = _T_262 ? medeleg : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_335 = _T_334 | _T_299; // @[Mux.scala 27:72]
  wire  _T_263 = 12'h105 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_300 = _T_263 ? stvec : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_336 = _T_335 | _T_300; // @[Mux.scala 27:72]
  wire  _T_264 = 12'h141 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_301 = _T_264 ? sepc : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_337 = _T_336 | _T_301; // @[Mux.scala 27:72]
  wire  _T_265 = 12'h342 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_302 = _T_265 ? mcause : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_338 = _T_337 | _T_302; // @[Mux.scala 27:72]
  wire  _T_266 = 12'h306 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_303 = _T_266 ? mcounteren : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_339 = _T_338 | _T_303; // @[Mux.scala 27:72]
  wire  _T_267 = 12'hf11 == addr; // @[LookupTree.scala 24:34]
  wire  _T_268 = 12'h104 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_231 = mie & sieMask; // @[RegMap.scala 48:84]
  wire [63:0] _T_305 = _T_268 ? _T_231 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_341 = _T_339 | _T_305; // @[Mux.scala 27:72]
  wire  _T_269 = 12'h144 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _GEN_79 = {{52'd0}, _T_113}; // @[RegMap.scala 48:84]
  wire [63:0] _T_232 = _GEN_79 & sieMask; // @[RegMap.scala 48:84]
  wire [63:0] _T_306 = _T_269 ? _T_232 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_342 = _T_341 | _T_306; // @[Mux.scala 27:72]
  wire  _T_270 = 12'h100 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_233 = mstatus & 64'h80000003000de122; // @[RegMap.scala 48:84]
  wire [63:0] _T_307 = _T_270 ? _T_233 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_343 = _T_342 | _T_307; // @[Mux.scala 27:72]
  wire  _T_271 = 12'h305 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_308 = _T_271 ? mtvec : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_344 = _T_343 | _T_308; // @[Mux.scala 27:72]
  wire  _T_272 = 12'h304 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_309 = _T_272 ? mie : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_345 = _T_344 | _T_309; // @[Mux.scala 27:72]
  wire  _T_273 = 12'hb01 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_310 = _T_273 ? perfCnts_1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_346 = _T_345 | _T_310; // @[Mux.scala 27:72]
  wire  _T_274 = 12'h3b3 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_311 = _T_274 ? pmpaddr3 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_347 = _T_346 | _T_311; // @[Mux.scala 27:72]
  wire  _T_275 = 12'h143 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_312 = _T_275 ? stval : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_348 = _T_347 | _T_312; // @[Mux.scala 27:72]
  wire  _T_276 = 12'h301 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_313 = _T_276 ? misa : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_349 = _T_348 | _T_313; // @[Mux.scala 27:72]
  wire  _T_277 = 12'h300 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_314 = _T_277 ? mstatus : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_350 = _T_349 | _T_314; // @[Mux.scala 27:72]
  wire  _T_278 = 12'hb00 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_315 = _T_278 ? perfCnts_0 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_351 = _T_350 | _T_315; // @[Mux.scala 27:72]
  wire  _T_279 = 12'h3b0 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_316 = _T_279 ? pmpaddr0 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_352 = _T_351 | _T_316; // @[Mux.scala 27:72]
  wire  _T_280 = 12'h344 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_317 = _T_280 ? _GEN_79 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_353 = _T_352 | _T_317; // @[Mux.scala 27:72]
  wire  _T_281 = 12'hb02 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_318 = _T_281 ? perfCnts_2 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_354 = _T_353 | _T_318; // @[Mux.scala 27:72]
  wire  _T_282 = 12'h3a3 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_319 = _T_282 ? pmpcfg3 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_355 = _T_354 | _T_319; // @[Mux.scala 27:72]
  wire  _T_283 = 12'h303 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_320 = _T_283 ? mideleg : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_356 = _T_355 | _T_320; // @[Mux.scala 27:72]
  wire  _T_284 = 12'h3b2 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_321 = _T_284 ? pmpaddr2 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_357 = _T_356 | _T_321; // @[Mux.scala 27:72]
  wire  _T_285 = 12'hf13 == addr; // @[LookupTree.scala 24:34]
  wire  _T_286 = 12'h3a1 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_323 = _T_286 ? pmpcfg1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_359 = _T_357 | _T_323; // @[Mux.scala 27:72]
  wire  _T_287 = 12'h340 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_324 = _T_287 ? mscratch : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_360 = _T_359 | _T_324; // @[Mux.scala 27:72]
  wire  _T_288 = 12'hf14 == addr; // @[LookupTree.scala 24:34]
  wire  _T_289 = 12'h341 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_326 = _T_289 ? mepc : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_362 = _T_360 | _T_326; // @[Mux.scala 27:72]
  wire  _T_290 = 12'h343 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_327 = _T_290 ? mtval : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_363 = _T_362 | _T_327; // @[Mux.scala 27:72]
  wire  _T_291 = 12'h106 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_328 = _T_291 ? scounteren : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_364 = _T_363 | _T_328; // @[Mux.scala 27:72]
  wire  _T_292 = 12'h3a0 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_329 = _T_292 ? pmpcfg0 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_365 = _T_364 | _T_329; // @[Mux.scala 27:72]
  wire  _T_293 = 12'h142 == addr; // @[LookupTree.scala 24:34]
  wire [63:0] _T_330 = _T_293 ? scause : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] rdata = _T_365 | _T_330; // @[Mux.scala 27:72]
  wire [63:0] _T_168 = rdata | io_in_bits_src1; // @[CSR.scala 460:30]
  wire [63:0] _T_169 = ~io_in_bits_src1; // @[CSR.scala 461:32]
  wire [63:0] _T_170 = rdata & _T_169; // @[CSR.scala 461:30]
  wire [63:0] _T_171 = rdata | csri; // @[CSR.scala 463:30]
  wire [63:0] _T_172 = ~csri; // @[CSR.scala 464:32]
  wire [63:0] _T_173 = rdata & _T_172; // @[CSR.scala 464:30]
  wire  _T_174 = 7'h1 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_175 = 7'h2 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_176 = 7'h3 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_177 = 7'h5 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_178 = 7'h6 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire  _T_179 = 7'h7 == io_in_bits_func; // @[LookupTree.scala 24:34]
  wire [63:0] _T_180 = _T_174 ? io_in_bits_src1 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_181 = _T_175 ? _T_168 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_182 = _T_176 ? _T_170 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_183 = _T_177 ? csri : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_184 = _T_178 ? _T_171 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_185 = _T_179 ? _T_173 : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_186 = _T_180 | _T_181; // @[Mux.scala 27:72]
  wire [63:0] _T_187 = _T_186 | _T_182; // @[Mux.scala 27:72]
  wire [63:0] _T_188 = _T_187 | _T_183; // @[Mux.scala 27:72]
  wire [63:0] _T_189 = _T_188 | _T_184; // @[Mux.scala 27:72]
  wire [63:0] wdata = _T_189 | _T_185; // @[Mux.scala 27:72]
  wire  _T_196 = wdata[63:60] == 4'h0; // @[CSR.scala 468:60]
  wire  _T_202 = wdata[63:60] == 4'h8; // @[CSR.scala 468:109]
  wire  satpLegalMode = _T_196 | _T_202; // @[CSR.scala 468:69]
  wire  _T_203 = io_in_bits_func != 7'h0; // @[CSR.scala 471:28]
  wire  _T_204 = io_in_valid & _T_203; // @[CSR.scala 471:20]
  wire  _T_205 = addr != 12'h180; // @[CSR.scala 471:56]
  wire  _T_206 = _T_205 | satpLegalMode; // @[CSR.scala 471:67]
  wire  wen = _T_204 & _T_206; // @[CSR.scala 471:47]
  wire  isIllegalMode = priviledgeMode < addr[9:8]; // @[CSR.scala 472:39]
  wire  _T_210 = io_in_bits_func == 7'h2; // @[CSR.scala 473:24]
  wire  _T_211 = io_in_bits_func == 7'h6; // @[CSR.scala 473:50]
  wire  _T_212 = _T_210 | _T_211; // @[CSR.scala 473:42]
  wire  _T_213 = io_in_bits_src1 == 64'h0; // @[CSR.scala 473:78]
  wire  justRead = _T_212 & _T_213; // @[CSR.scala 473:70]
  wire  _T_215 = addr[11:10] == 2'h3; // @[CSR.scala 474:45]
  wire  _T_216 = wen & _T_215; // @[CSR.scala 474:28]
  wire  _T_217 = ~justRead; // @[CSR.scala 474:61]
  wire  isIllegalWrite = _T_216 & _T_217; // @[CSR.scala 474:58]
  wire  isIllegalAccess = isIllegalMode | isIllegalWrite; // @[CSR.scala 475:39]
  wire  _T_218 = ~isIllegalAccess; // @[CSR.scala 477:54]
  wire  _T_219 = wen & _T_218; // @[CSR.scala 477:51]
  wire  _T_368 = addr == 12'h180; // @[RegMap.scala 50:65]
  wire  _T_369 = _T_219 & _T_368; // @[RegMap.scala 50:56]
  wire  _T_374 = addr == 12'h3b1; // @[RegMap.scala 50:65]
  wire  _T_375 = _T_219 & _T_374; // @[RegMap.scala 50:56]
  wire  _T_380 = addr == 12'h3a2; // @[RegMap.scala 50:65]
  wire  _T_381 = _T_219 & _T_380; // @[RegMap.scala 50:56]
  wire  _T_386 = addr == 12'h140; // @[RegMap.scala 50:65]
  wire  _T_387 = _T_219 & _T_386; // @[RegMap.scala 50:56]
  wire  _T_392 = addr == 12'h302; // @[RegMap.scala 50:65]
  wire  _T_393 = _T_219 & _T_392; // @[RegMap.scala 50:56]
  wire [63:0] _T_394 = wdata & 64'hbbff; // @[BitUtils.scala 32:13]
  wire [63:0] _T_396 = medeleg & 64'h4400; // @[BitUtils.scala 32:36]
  wire [63:0] _T_397 = _T_394 | _T_396; // @[BitUtils.scala 32:25]
  wire  _T_398 = addr == 12'h105; // @[RegMap.scala 50:65]
  wire  _T_399 = _T_219 & _T_398; // @[RegMap.scala 50:56]
  wire  _T_404 = addr == 12'h141; // @[RegMap.scala 50:65]
  wire  _T_405 = _T_219 & _T_404; // @[RegMap.scala 50:56]
  wire  _T_410 = addr == 12'h342; // @[RegMap.scala 50:65]
  wire  _T_411 = _T_219 & _T_410; // @[RegMap.scala 50:56]
  wire  _T_416 = addr == 12'h306; // @[RegMap.scala 50:65]
  wire  _T_417 = _T_219 & _T_416; // @[RegMap.scala 50:56]
  wire  _T_422 = addr == 12'h104; // @[RegMap.scala 50:65]
  wire  _T_423 = _T_219 & _T_422; // @[RegMap.scala 50:56]
  wire [63:0] _T_424 = wdata & sieMask; // @[BitUtils.scala 32:13]
  wire [63:0] _T_425 = ~sieMask; // @[BitUtils.scala 32:38]
  wire [63:0] _T_426 = mie & _T_425; // @[BitUtils.scala 32:36]
  wire [63:0] _T_427 = _T_424 | _T_426; // @[BitUtils.scala 32:25]
  wire  _T_428 = addr == 12'h100; // @[RegMap.scala 50:65]
  wire  _T_429 = _T_219 & _T_428; // @[RegMap.scala 50:56]
  wire [63:0] _T_430 = wdata & 64'hc6122; // @[BitUtils.scala 32:13]
  wire [63:0] _T_432 = mstatus & 64'h39edd; // @[BitUtils.scala 32:36]
  wire [63:0] _T_433 = _T_430 | _T_432; // @[BitUtils.scala 32:25]
  wire  _T_461 = _T_433[14:13] == 2'h3; // @[CSR.scala 301:40]
  wire [63:0] _T_463 = {_T_461,_T_433[62:0]}; // @[Cat.scala 29:58]
  wire  _T_464 = addr == 12'h305; // @[RegMap.scala 50:65]
  wire  _T_465 = _T_219 & _T_464; // @[RegMap.scala 50:56]
  wire  _T_470 = addr == 12'h304; // @[RegMap.scala 50:65]
  wire  _T_471 = _T_219 & _T_470; // @[RegMap.scala 50:56]
  wire  _T_476 = addr == 12'hb01; // @[RegMap.scala 50:65]
  wire  _T_477 = _T_219 & _T_476; // @[RegMap.scala 50:56]
  wire  _T_482 = addr == 12'h3b3; // @[RegMap.scala 50:65]
  wire  _T_483 = _T_219 & _T_482; // @[RegMap.scala 50:56]
  wire  _T_488 = addr == 12'h143; // @[RegMap.scala 50:65]
  wire  _T_489 = _T_219 & _T_488; // @[RegMap.scala 50:56]
  wire [63:0] _GEN_17 = _T_489 ? wdata : stval; // @[RegMap.scala 50:72]
  wire  _T_494 = addr == 12'h301; // @[RegMap.scala 50:65]
  wire  _T_495 = _T_219 & _T_494; // @[RegMap.scala 50:56]
  wire  _T_500 = addr == 12'h300; // @[RegMap.scala 50:65]
  wire  _T_501 = _T_219 & _T_500; // @[RegMap.scala 50:56]
  wire  _T_533 = wdata[14:13] == 2'h3; // @[CSR.scala 301:40]
  wire [63:0] _T_535 = {_T_533,wdata[62:0]}; // @[Cat.scala 29:58]
  wire  _T_542 = addr == 12'h3b0; // @[RegMap.scala 50:65]
  wire  _T_543 = _T_219 & _T_542; // @[RegMap.scala 50:56]
  wire  _T_548 = addr == 12'hb02; // @[RegMap.scala 50:65]
  wire  _T_549 = _T_219 & _T_548; // @[RegMap.scala 50:56]
  wire  _T_554 = addr == 12'h3a3; // @[RegMap.scala 50:65]
  wire  _T_555 = _T_219 & _T_554; // @[RegMap.scala 50:56]
  wire  _T_560 = addr == 12'h303; // @[RegMap.scala 50:65]
  wire  _T_561 = _T_219 & _T_560; // @[RegMap.scala 50:56]
  wire [63:0] _T_562 = wdata & 64'h222; // @[BitUtils.scala 32:13]
  wire [63:0] _T_564 = mideleg & 64'h1dd; // @[BitUtils.scala 32:36]
  wire [63:0] _T_565 = _T_562 | _T_564; // @[BitUtils.scala 32:25]
  wire  _T_566 = addr == 12'h3b2; // @[RegMap.scala 50:65]
  wire  _T_567 = _T_219 & _T_566; // @[RegMap.scala 50:56]
  wire  _T_572 = addr == 12'h3a1; // @[RegMap.scala 50:65]
  wire  _T_573 = _T_219 & _T_572; // @[RegMap.scala 50:56]
  wire  _T_578 = addr == 12'h340; // @[RegMap.scala 50:65]
  wire  _T_579 = _T_219 & _T_578; // @[RegMap.scala 50:56]
  wire  _T_584 = addr == 12'h341; // @[RegMap.scala 50:65]
  wire  _T_585 = _T_219 & _T_584; // @[RegMap.scala 50:56]
  wire  _T_590 = addr == 12'h343; // @[RegMap.scala 50:65]
  wire  _T_591 = _T_219 & _T_590; // @[RegMap.scala 50:56]
  wire [63:0] _GEN_29 = _T_591 ? wdata : mtval; // @[RegMap.scala 50:72]
  wire  _T_596 = addr == 12'h106; // @[RegMap.scala 50:65]
  wire  _T_597 = _T_219 & _T_596; // @[RegMap.scala 50:56]
  wire  _T_602 = addr == 12'h3a0; // @[RegMap.scala 50:65]
  wire  _T_603 = _T_219 & _T_602; // @[RegMap.scala 50:56]
  wire  _T_608 = addr == 12'h142; // @[RegMap.scala 50:65]
  wire  _T_609 = _T_219 & _T_608; // @[RegMap.scala 50:56]
  wire  _T_615 = _T_257 ? 1'h0 : 1'h1; // @[Mux.scala 80:57]
  wire  _T_617 = _T_258 ? 1'h0 : _T_615; // @[Mux.scala 80:57]
  wire  _T_619 = _T_259 ? 1'h0 : _T_617; // @[Mux.scala 80:57]
  wire  _T_621 = _T_260 ? 1'h0 : _T_619; // @[Mux.scala 80:57]
  wire  _T_623 = _T_261 ? 1'h0 : _T_621; // @[Mux.scala 80:57]
  wire  _T_625 = _T_262 ? 1'h0 : _T_623; // @[Mux.scala 80:57]
  wire  _T_627 = _T_263 ? 1'h0 : _T_625; // @[Mux.scala 80:57]
  wire  _T_629 = _T_264 ? 1'h0 : _T_627; // @[Mux.scala 80:57]
  wire  _T_631 = _T_265 ? 1'h0 : _T_629; // @[Mux.scala 80:57]
  wire  _T_633 = _T_266 ? 1'h0 : _T_631; // @[Mux.scala 80:57]
  wire  _T_635 = _T_267 ? 1'h0 : _T_633; // @[Mux.scala 80:57]
  wire  _T_637 = _T_268 ? 1'h0 : _T_635; // @[Mux.scala 80:57]
  wire  _T_639 = _T_269 ? 1'h0 : _T_637; // @[Mux.scala 80:57]
  wire  _T_641 = _T_270 ? 1'h0 : _T_639; // @[Mux.scala 80:57]
  wire  _T_643 = _T_271 ? 1'h0 : _T_641; // @[Mux.scala 80:57]
  wire  _T_645 = _T_272 ? 1'h0 : _T_643; // @[Mux.scala 80:57]
  wire  _T_647 = _T_273 ? 1'h0 : _T_645; // @[Mux.scala 80:57]
  wire  _T_649 = _T_274 ? 1'h0 : _T_647; // @[Mux.scala 80:57]
  wire  _T_651 = _T_275 ? 1'h0 : _T_649; // @[Mux.scala 80:57]
  wire  _T_653 = _T_276 ? 1'h0 : _T_651; // @[Mux.scala 80:57]
  wire  _T_655 = _T_277 ? 1'h0 : _T_653; // @[Mux.scala 80:57]
  wire  _T_657 = _T_278 ? 1'h0 : _T_655; // @[Mux.scala 80:57]
  wire  _T_659 = _T_279 ? 1'h0 : _T_657; // @[Mux.scala 80:57]
  wire  _T_661 = _T_280 ? 1'h0 : _T_659; // @[Mux.scala 80:57]
  wire  _T_663 = _T_281 ? 1'h0 : _T_661; // @[Mux.scala 80:57]
  wire  _T_665 = _T_282 ? 1'h0 : _T_663; // @[Mux.scala 80:57]
  wire  _T_667 = _T_283 ? 1'h0 : _T_665; // @[Mux.scala 80:57]
  wire  _T_669 = _T_284 ? 1'h0 : _T_667; // @[Mux.scala 80:57]
  wire  _T_671 = _T_285 ? 1'h0 : _T_669; // @[Mux.scala 80:57]
  wire  _T_673 = _T_286 ? 1'h0 : _T_671; // @[Mux.scala 80:57]
  wire  _T_675 = _T_287 ? 1'h0 : _T_673; // @[Mux.scala 80:57]
  wire  _T_677 = _T_288 ? 1'h0 : _T_675; // @[Mux.scala 80:57]
  wire  _T_679 = _T_289 ? 1'h0 : _T_677; // @[Mux.scala 80:57]
  wire  _T_681 = _T_290 ? 1'h0 : _T_679; // @[Mux.scala 80:57]
  wire  _T_683 = _T_291 ? 1'h0 : _T_681; // @[Mux.scala 80:57]
  wire  _T_685 = _T_292 ? 1'h0 : _T_683; // @[Mux.scala 80:57]
  wire  isIllegalAddr = _T_293 ? 1'h0 : _T_685; // @[Mux.scala 80:57]
  wire  resetSatp = _T_368 & wen; // @[CSR.scala 479:35]
  wire  _T_700 = addr == 12'h344; // @[RegMap.scala 50:65]
  wire  _T_701 = _T_219 & _T_700; // @[RegMap.scala 50:56]
  wire [63:0] _T_702 = wdata & 64'h77f; // @[BitUtils.scala 32:13]
  wire [63:0] _T_704 = mipReg & 64'h80; // @[BitUtils.scala 32:36]
  wire [63:0] _T_705 = _T_702 | _T_704; // @[BitUtils.scala 32:25]
  wire  _T_706 = addr == 12'h144; // @[RegMap.scala 50:65]
  wire  _T_707 = _T_219 & _T_706; // @[RegMap.scala 50:56]
  wire [63:0] _T_710 = mipReg & _T_425; // @[BitUtils.scala 32:36]
  wire [63:0] _T_711 = _T_424 | _T_710; // @[BitUtils.scala 32:25]
  wire  _T_712 = addr == 12'h1; // @[CSR.scala 492:23]
  wire  _T_713 = io_in_bits_func == 7'h0; // @[CSR.scala 492:46]
  wire  isEbreak = _T_712 & _T_713; // @[CSR.scala 492:38]
  wire  _T_716 = addr == 12'h0; // @[CSR.scala 493:22]
  wire  isEcall = _T_716 & _T_713; // @[CSR.scala 493:36]
  wire  isMret = _T_392 & _T_713; // @[CSR.scala 494:36]
  wire  _T_724 = addr == 12'h102; // @[CSR.scala 495:21]
  wire  isSret = _T_724 & _T_713; // @[CSR.scala 495:36]
  wire  _T_728 = addr == 12'h2; // @[CSR.scala 496:21]
  wire  isUret = _T_728 & _T_713; // @[CSR.scala 496:36]
  wire  hasInstrPageFault = io_cfIn_exceptionVec_12 & io_in_valid; // @[CSR.scala 553:63]
  wire  _T_759 = hasInstrPageFault | io_dmemMMU_loadPF; // @[CSR.scala 562:26]
  wire  _T_760 = _T_759 | io_dmemMMU_storePF; // @[CSR.scala 562:46]
  wire [38:0] _T_762 = io_cfIn_pc + 39'h2; // @[CSR.scala 563:88]
  wire [24:0] _T_766 = _T_762[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_767 = {_T_766,_T_762}; // @[Cat.scala 29:58]
  wire [24:0] _T_771 = io_cfIn_pc[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_772 = {_T_771,io_cfIn_pc}; // @[Cat.scala 29:58]
  wire [63:0] _T_773 = io_cfIn_crossPageIPFFix ? _T_767 : _T_772; // @[CSR.scala 563:42]
  wire [24:0] _T_776 = io_dmemMMU_addr[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_777 = {_T_776,io_dmemMMU_addr}; // @[Cat.scala 29:58]
  wire [63:0] _T_778 = hasInstrPageFault ? _T_773 : _T_777; // @[CSR.scala 563:19]
  wire  _T_779 = priviledgeMode == 2'h3; // @[CSR.scala 564:25]
  wire  _T_796 = io_cfIn_exceptionVec_4 | io_cfIn_exceptionVec_6; // @[CSR.scala 572:30]
  wire [38:0] dmemAddrMisalignedAddr = LSUADDR[38:0]; // @[CSR.scala 541:36 CSR.scala 559:28]
  wire [24:0] _T_799 = dmemAddrMisalignedAddr[38] ? 25'h1ffffff : 25'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_800 = {_T_799,dmemAddrMisalignedAddr}; // @[Cat.scala 29:58]
  wire  mipRaiseIntr_e_s = mip_e_s | meip_0; // @[CSR.scala 596:31]
  wire [11:0] _T_828 = {mip_e_m,mip_e_h,mipRaiseIntr_e_s,mip_e_u,mip_t_m,mip_t_h,_T_107}; // @[CSR.scala 598:41]
  wire [63:0] _GEN_80 = {{52'd0}, _T_828}; // @[CSR.scala 598:26]
  wire [63:0] ideleg = mideleg & _GEN_80; // @[CSR.scala 598:26]
  wire  _T_893 = priviledgeMode == 2'h1; // @[CSR.scala 599:72]
  wire  _T_894 = _T_893 & mstatusStruct_ie_s; // @[CSR.scala 599:83]
  wire  _T_895 = priviledgeMode < 2'h1; // @[CSR.scala 599:125]
  wire  _T_896 = _T_894 | _T_895; // @[CSR.scala 599:106]
  wire  _T_898 = _T_779 & mstatusStruct_ie_m; // @[CSR.scala 600:64]
  wire  _T_899 = priviledgeMode < 2'h3; // @[CSR.scala 600:106]
  wire  _T_900 = _T_898 | _T_899; // @[CSR.scala 600:87]
  wire  intrVecEnable_0 = ideleg[0] ? _T_896 : _T_900; // @[CSR.scala 599:51]
  wire  intrVecEnable_1 = ideleg[1] ? _T_896 : _T_900; // @[CSR.scala 599:51]
  wire  intrVecEnable_2 = ideleg[2] ? _T_896 : _T_900; // @[CSR.scala 599:51]
  wire  intrVecEnable_3 = ideleg[3] ? _T_896 : _T_900; // @[CSR.scala 599:51]
  wire  intrVecEnable_4 = ideleg[4] ? _T_896 : _T_900; // @[CSR.scala 599:51]
  wire  intrVecEnable_5 = ideleg[5] ? _T_896 : _T_900; // @[CSR.scala 599:51]
  wire  intrVecEnable_6 = ideleg[6] ? _T_896 : _T_900; // @[CSR.scala 599:51]
  wire  intrVecEnable_7 = ideleg[7] ? _T_896 : _T_900; // @[CSR.scala 599:51]
  wire  intrVecEnable_8 = ideleg[8] ? _T_896 : _T_900; // @[CSR.scala 599:51]
  wire  intrVecEnable_9 = ideleg[9] ? _T_896 : _T_900; // @[CSR.scala 599:51]
  wire  intrVecEnable_10 = ideleg[10] ? _T_896 : _T_900; // @[CSR.scala 599:51]
  wire  intrVecEnable_11 = ideleg[11] ? _T_896 : _T_900; // @[CSR.scala 599:51]
  wire [11:0] _T_1013 = mie[11:0] & _T_828; // @[CSR.scala 604:27]
  wire [5:0] _T_1018 = {intrVecEnable_5,intrVecEnable_4,intrVecEnable_3,intrVecEnable_2,intrVecEnable_1,intrVecEnable_0}; // @[CSR.scala 604:65]
  wire [11:0] _T_1024 = {intrVecEnable_11,intrVecEnable_10,intrVecEnable_9,intrVecEnable_8,intrVecEnable_7,intrVecEnable_6,_T_1018}; // @[CSR.scala 604:65]
  wire [11:0] intrVec = _T_1013 & _T_1024; // @[CSR.scala 604:49]
  wire [2:0] _T_1025 = io_cfIn_intrVec_4 ? 3'h4 : 3'h0; // @[CSR.scala 608:69]
  wire [3:0] _T_1026 = io_cfIn_intrVec_8 ? 4'h8 : {{1'd0}, _T_1025}; // @[CSR.scala 608:69]
  wire [3:0] _T_1027 = io_cfIn_intrVec_0 ? 4'h0 : _T_1026; // @[CSR.scala 608:69]
  wire [3:0] _T_1028 = io_cfIn_intrVec_5 ? 4'h5 : _T_1027; // @[CSR.scala 608:69]
  wire [3:0] _T_1029 = io_cfIn_intrVec_9 ? 4'h9 : _T_1028; // @[CSR.scala 608:69]
  wire [3:0] _T_1030 = io_cfIn_intrVec_1 ? 4'h1 : _T_1029; // @[CSR.scala 608:69]
  wire [3:0] _T_1031 = io_cfIn_intrVec_7 ? 4'h7 : _T_1030; // @[CSR.scala 608:69]
  wire [3:0] _T_1032 = io_cfIn_intrVec_11 ? 4'hb : _T_1031; // @[CSR.scala 608:69]
  wire [3:0] intrNO = io_cfIn_intrVec_3 ? 4'h3 : _T_1032; // @[CSR.scala 608:69]
  wire [5:0] _T_1037 = {io_cfIn_intrVec_5,io_cfIn_intrVec_4,io_cfIn_intrVec_3,io_cfIn_intrVec_2,io_cfIn_intrVec_1,io_cfIn_intrVec_0}; // @[CSR.scala 610:35]
  wire [11:0] _T_1043 = {io_cfIn_intrVec_11,io_cfIn_intrVec_10,io_cfIn_intrVec_9,io_cfIn_intrVec_8,io_cfIn_intrVec_7,io_cfIn_intrVec_6,_T_1037}; // @[CSR.scala 610:35]
  wire  raiseIntr = |_T_1043; // @[CSR.scala 610:42]
  wire  csrExceptionVec_3 = io_in_valid & isEbreak; // @[CSR.scala 617:46]
  wire  _T_1046 = _T_779 & io_in_valid; // @[CSR.scala 618:55]
  wire  csrExceptionVec_11 = _T_1046 & isEcall; // @[CSR.scala 618:70]
  wire  _T_1049 = _T_893 & io_in_valid; // @[CSR.scala 619:55]
  wire  csrExceptionVec_9 = _T_1049 & isEcall; // @[CSR.scala 619:70]
  wire  _T_1051 = priviledgeMode == 2'h0; // @[CSR.scala 620:45]
  wire  _T_1052 = _T_1051 & io_in_valid; // @[CSR.scala 620:55]
  wire  csrExceptionVec_8 = _T_1052 & isEcall; // @[CSR.scala 620:70]
  wire  _T_1054 = isIllegalAddr | isIllegalAccess; // @[CSR.scala 621:51]
  wire  csrExceptionVec_2 = _T_1054 & wen; // @[CSR.scala 621:71]
  wire [7:0] _T_1064 = {4'h0,csrExceptionVec_3,csrExceptionVec_2,2'h0}; // @[CSR.scala 625:49]
  wire [15:0] _T_1072 = {io_dmemMMU_storePF,1'h0,io_dmemMMU_loadPF,1'h0,csrExceptionVec_11,1'h0,csrExceptionVec_9,csrExceptionVec_8,_T_1064}; // @[CSR.scala 625:49]
  wire [7:0] _T_1079 = {1'h0,io_cfIn_exceptionVec_6,1'h0,io_cfIn_exceptionVec_4,1'h0,io_cfIn_exceptionVec_2,io_cfIn_exceptionVec_1,1'h0}; // @[CSR.scala 625:76]
  wire [15:0] _T_1087 = {2'h0,1'h0,io_cfIn_exceptionVec_12,4'h0,_T_1079}; // @[CSR.scala 625:76]
  wire [15:0] raiseExceptionVec = _T_1072 | _T_1087; // @[CSR.scala 625:52]
  wire  raiseException = |raiseExceptionVec; // @[CSR.scala 626:42]
  wire [2:0] _T_1089 = raiseExceptionVec[5] ? 3'h5 : 3'h0; // @[CSR.scala 627:74]
  wire [2:0] _T_1091 = raiseExceptionVec[7] ? 3'h7 : _T_1089; // @[CSR.scala 627:74]
  wire [3:0] _T_1093 = raiseExceptionVec[13] ? 4'hd : {{1'd0}, _T_1091}; // @[CSR.scala 627:74]
  wire [3:0] _T_1095 = raiseExceptionVec[15] ? 4'hf : _T_1093; // @[CSR.scala 627:74]
  wire [3:0] _T_1097 = raiseExceptionVec[4] ? 4'h4 : _T_1095; // @[CSR.scala 627:74]
  wire [3:0] _T_1099 = raiseExceptionVec[6] ? 4'h6 : _T_1097; // @[CSR.scala 627:74]
  wire [3:0] _T_1101 = raiseExceptionVec[8] ? 4'h8 : _T_1099; // @[CSR.scala 627:74]
  wire [3:0] _T_1103 = raiseExceptionVec[9] ? 4'h9 : _T_1101; // @[CSR.scala 627:74]
  wire [3:0] _T_1105 = raiseExceptionVec[11] ? 4'hb : _T_1103; // @[CSR.scala 627:74]
  wire [3:0] _T_1107 = raiseExceptionVec[0] ? 4'h0 : _T_1105; // @[CSR.scala 627:74]
  wire [3:0] _T_1109 = raiseExceptionVec[2] ? 4'h2 : _T_1107; // @[CSR.scala 627:74]
  wire [3:0] _T_1111 = raiseExceptionVec[1] ? 4'h1 : _T_1109; // @[CSR.scala 627:74]
  wire [3:0] _T_1113 = raiseExceptionVec[12] ? 4'hc : _T_1111; // @[CSR.scala 627:74]
  wire [3:0] exceptionNO = raiseExceptionVec[3] ? 4'h3 : _T_1113; // @[CSR.scala 627:74]
  wire [63:0] _T_1115 = {raiseIntr, 63'h0}; // @[CSR.scala 630:28]
  wire [3:0] _T_1116 = raiseIntr ? intrNO : exceptionNO; // @[CSR.scala 630:46]
  wire [63:0] _GEN_81 = {{60'd0}, _T_1116}; // @[CSR.scala 630:41]
  wire [63:0] causeNO = _T_1115 | _GEN_81; // @[CSR.scala 630:41]
  wire  _T_1118 = raiseException | raiseIntr; // @[CSR.scala 633:44]
  wire  raiseExceptionIntr = _T_1118 & io_instrValid; // @[CSR.scala 633:58]
  wire  _T_1120 = io_in_valid & _T_713; // @[CSR.scala 636:31]
  wire  _T_1121 = _T_1120 | raiseExceptionIntr; // @[CSR.scala 636:58]
  wire [38:0] _T_1124 = io_cfIn_pc + 39'h4; // @[CSR.scala 638:51]
  wire [63:0] deleg = raiseIntr ? mideleg : medeleg; // @[CSR.scala 648:18]
  wire [63:0] _T_1217 = deleg >> causeNO[3:0]; // @[CSR.scala 650:22]
  wire  delegS = _T_1217[0] & _T_899; // @[CSR.scala 650:38]
  wire [63:0] _T_1227 = delegS ? stvec : mtvec; // @[CSR.scala 654:20]
  wire [38:0] trapTarget = _T_1227[38:0]; // @[CSR.scala 654:42]
  wire  _T_1388 = io_in_valid & isUret; // @[CSR.scala 685:15]
  wire  _T_1308 = io_in_valid & isSret; // @[CSR.scala 672:15]
  wire  _T_1229 = io_in_valid & isMret; // @[CSR.scala 659:15]
  wire [38:0] _GEN_47 = _T_1308 ? sepc[38:0] : mepc[38:0]; // @[CSR.scala 672:26]
  wire [38:0] retTarget = _T_1388 ? 39'h0 : _GEN_47; // @[CSR.scala 685:26]
  wire [38:0] _T_1125 = raiseExceptionIntr ? trapTarget : retTarget; // @[CSR.scala 638:61]
  wire  _T_1222 = _T_760 | io_cfIn_exceptionVec_4; // @[CSR.scala 651:78]
  wire  _T_1223 = _T_1222 | io_cfIn_exceptionVec_6; // @[CSR.scala 651:103]
  wire  _T_1224 = ~_T_1223; // @[CSR.scala 651:17]
  wire  tvalWen = _T_1224 | raiseIntr; // @[CSR.scala 651:130]
  wire [5:0] _T_1288 = {mstatusStruct_pie_s,mstatusStruct_pie_u,mstatusStruct_pie_m,mstatusStruct_ie_h,mstatusStruct_ie_s,mstatusStruct_ie_u}; // @[CSR.scala 667:27]
  wire [14:0] _T_1294 = {mstatusStruct_fs,2'h0,mstatusStruct_hpp,mstatusStruct_spp,1'h1,mstatusStruct_pie_h,_T_1288}; // @[CSR.scala 667:27]
  wire [6:0] _T_1299 = {mstatusStruct_tw,mstatusStruct_tvm,mstatusStruct_mxr,mstatusStruct_sum,mstatusStruct_mprv,mstatusStruct_xs}; // @[CSR.scala 667:27]
  wire [63:0] _T_1306 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,mstatusStruct_pad0,mstatusStruct_tsr,_T_1299,_T_1294}; // @[CSR.scala 667:27]
  wire [1:0] _T_1363 = {1'h0,mstatusStruct_spp}; // @[Cat.scala 29:58]
  wire [5:0] _T_1368 = {1'h1,mstatusStruct_pie_u,mstatusStruct_ie_m,mstatusStruct_ie_h,mstatusStruct_pie_s,mstatusStruct_ie_u}; // @[CSR.scala 680:27]
  wire [14:0] _T_1374 = {mstatusStruct_fs,mstatusStruct_mpp,mstatusStruct_hpp,1'h0,mstatusStruct_pie_m,mstatusStruct_pie_h,_T_1368}; // @[CSR.scala 680:27]
  wire [63:0] _T_1386 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,mstatusStruct_pad0,mstatusStruct_tsr,_T_1299,_T_1374}; // @[CSR.scala 680:27]
  wire [5:0] _T_1447 = {mstatusStruct_pie_s,1'h1,mstatusStruct_ie_m,mstatusStruct_ie_h,mstatusStruct_ie_s,mstatusStruct_pie_u}; // @[CSR.scala 692:27]
  wire [14:0] _T_1453 = {mstatusStruct_fs,mstatusStruct_mpp,mstatusStruct_hpp,mstatusStruct_spp,mstatusStruct_pie_m,mstatusStruct_pie_h,_T_1447}; // @[CSR.scala 692:27]
  wire [63:0] _T_1465 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,mstatusStruct_pad0,mstatusStruct_tsr,_T_1299,_T_1453}; // @[CSR.scala 692:27]
  wire [1:0] _GEN_55 = delegS ? priviledgeMode : {{1'd0}, mstatusStruct_spp}; // @[CSR.scala 700:19]
  wire  _GEN_56 = delegS ? mstatusStruct_ie_s : mstatusStruct_pie_s; // @[CSR.scala 700:19]
  wire  _GEN_57 = delegS ? 1'h0 : mstatusStruct_ie_s; // @[CSR.scala 700:19]
  wire [1:0] _GEN_62 = delegS ? mstatusStruct_mpp : priviledgeMode; // @[CSR.scala 700:19]
  wire  _GEN_63 = delegS ? mstatusStruct_pie_m : mstatusStruct_ie_m; // @[CSR.scala 700:19]
  wire  _GEN_64 = delegS & mstatusStruct_ie_m; // @[CSR.scala 700:19]
  wire [5:0] _T_1533 = {_GEN_56,mstatusStruct_pie_u,_GEN_64,mstatusStruct_ie_h,_GEN_57,mstatusStruct_ie_u}; // @[CSR.scala 727:27]
  wire [14:0] _T_1539 = {mstatusStruct_fs,_GEN_62,mstatusStruct_hpp,_GEN_55[0],_GEN_63,mstatusStruct_pie_h,_T_1533}; // @[CSR.scala 727:27]
  wire [63:0] _T_1551 = {mstatusStruct_sd,mstatusStruct_pad1,mstatusStruct_sxl,mstatusStruct_uxl,mstatusStruct_pad0,mstatusStruct_tsr,_T_1299,_T_1539}; // @[CSR.scala 727:27]
  wire [63:0] _T_1553 = perfCnts_0 + 64'h1; // @[CSR.scala 836:71]
  wire  _T_1560 = 1'h1;
  wire [63:0] _T_1557 = perfCnts_2 + 64'h1; // @[CSR.scala 836:71]
  wire [63:0] _T_1559 = perfCnts_2 + 64'h2; // @[CSR.scala 844:86]
  assign io_out_valid = io_in_valid; // @[CSR.scala 731:16]
  assign io_out_bits = _T_365 | _T_330; // @[CSR.scala 480:15]
  assign io_redirect_target = resetSatp ? _T_1124 : _T_1125; // @[CSR.scala 638:22]
  assign io_redirect_valid = _T_1121 | resetSatp; // @[CSR.scala 636:21]
  assign io_imemMMU_priviledgeMode = priviledgeMode; // @[CSR.scala 527:29]
  assign io_dmemMMU_priviledgeMode = mstatusStruct_mprv ? mstatusStruct_mpp : priviledgeMode; // @[CSR.scala 528:29]
  assign io_dmemMMU_status_sum = mstatus[18]; // @[CSR.scala 530:25]
  assign io_dmemMMU_status_mxr = mstatus[19]; // @[CSR.scala 532:25]
  assign io_wenFix = |raiseExceptionVec; // @[CSR.scala 628:13]
  assign perfCnts_2_0 = perfCnts_2;
  assign satp_0 = satp;
  assign intrVec_0 = intrVec;
  assign lrAddr_0 = lrAddr;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  mtvec = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  mcounteren = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  mcause = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  mtval = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  mepc = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  mie = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mipReg = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  misa = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  mstatus = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  medeleg = _RAND_9[63:0];
  _RAND_10 = {2{`RANDOM}};
  mideleg = _RAND_10[63:0];
  _RAND_11 = {2{`RANDOM}};
  mscratch = _RAND_11[63:0];
  _RAND_12 = {2{`RANDOM}};
  pmpcfg0 = _RAND_12[63:0];
  _RAND_13 = {2{`RANDOM}};
  pmpcfg1 = _RAND_13[63:0];
  _RAND_14 = {2{`RANDOM}};
  pmpcfg2 = _RAND_14[63:0];
  _RAND_15 = {2{`RANDOM}};
  pmpcfg3 = _RAND_15[63:0];
  _RAND_16 = {2{`RANDOM}};
  pmpaddr0 = _RAND_16[63:0];
  _RAND_17 = {2{`RANDOM}};
  pmpaddr1 = _RAND_17[63:0];
  _RAND_18 = {2{`RANDOM}};
  pmpaddr2 = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  pmpaddr3 = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  stvec = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  satp = _RAND_21[63:0];
  _RAND_22 = {2{`RANDOM}};
  sepc = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  scause = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  stval = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  sscratch = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  scounteren = _RAND_26[63:0];
  _RAND_27 = {1{`RANDOM}};
  lr = _RAND_27[0:0];
  _RAND_28 = {2{`RANDOM}};
  lrAddr = _RAND_28[63:0];
  _RAND_29 = {1{`RANDOM}};
  priviledgeMode = _RAND_29[1:0];
  _RAND_30 = {2{`RANDOM}};
  perfCnts_0 = _RAND_30[63:0];
  _RAND_31 = {2{`RANDOM}};
  perfCnts_1 = _RAND_31[63:0];
  _RAND_32 = {2{`RANDOM}};
  perfCnts_2 = _RAND_32[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      mtvec <= 64'h0;
    end else if (_T_465) begin
      mtvec <= wdata;
    end
    if (reset) begin
      mcounteren <= 64'h0;
    end else if (_T_417) begin
      mcounteren <= wdata;
    end
    if (reset) begin
      mcause <= 64'h0;
    end else if (raiseExceptionIntr) begin
      if (delegS) begin
        if (_T_411) begin
          mcause <= wdata;
        end
      end else begin
        mcause <= causeNO;
      end
    end else if (_T_411) begin
      mcause <= wdata;
    end
    if (reset) begin
      mtval <= 64'h0;
    end else if (raiseExceptionIntr) begin
      if (delegS) begin
        if (_T_796) begin
          mtval <= _T_800;
        end else if (_T_760) begin
          if (_T_779) begin
            if (hasInstrPageFault) begin
              if (io_cfIn_crossPageIPFFix) begin
                mtval <= _T_767;
              end else begin
                mtval <= _T_772;
              end
            end else begin
              mtval <= _T_777;
            end
          end else if (_T_591) begin
            mtval <= wdata;
          end
        end else if (_T_591) begin
          mtval <= wdata;
        end
      end else if (tvalWen) begin
        mtval <= 64'h0;
      end else if (_T_796) begin
        mtval <= _T_800;
      end else if (_T_760) begin
        if (_T_779) begin
          if (hasInstrPageFault) begin
            if (io_cfIn_crossPageIPFFix) begin
              mtval <= _T_767;
            end else begin
              mtval <= _T_772;
            end
          end else begin
            mtval <= _T_777;
          end
        end else if (_T_591) begin
          mtval <= wdata;
        end
      end else if (_T_591) begin
        mtval <= wdata;
      end
    end else if (_T_796) begin
      mtval <= _T_800;
    end else if (_T_760) begin
      if (_T_779) begin
        if (hasInstrPageFault) begin
          if (io_cfIn_crossPageIPFFix) begin
            mtval <= _T_767;
          end else begin
            mtval <= _T_772;
          end
        end else begin
          mtval <= _T_777;
        end
      end else begin
        mtval <= _GEN_29;
      end
    end else begin
      mtval <= _GEN_29;
    end
    if (raiseExceptionIntr) begin
      if (delegS) begin
        if (_T_585) begin
          mepc <= wdata;
        end
      end else begin
        mepc <= _T_772;
      end
    end else if (_T_585) begin
      mepc <= wdata;
    end
    if (reset) begin
      mie <= 64'h0;
    end else if (_T_471) begin
      mie <= wdata;
    end else if (_T_423) begin
      mie <= _T_427;
    end
    if (reset) begin
      mipReg <= 64'h0;
    end else if (_T_707) begin
      mipReg <= _T_711;
    end else if (_T_701) begin
      mipReg <= _T_705;
    end
    if (reset) begin
      misa <= 64'h8000000000141105;
    end else if (_T_495) begin
      misa <= wdata;
    end
    if (reset) begin
      mstatus <= 64'h1800;
    end else if (raiseExceptionIntr) begin
      mstatus <= _T_1551;
    end else if (_T_1388) begin
      mstatus <= _T_1465;
    end else if (_T_1308) begin
      mstatus <= _T_1386;
    end else if (_T_1229) begin
      mstatus <= _T_1306;
    end else if (_T_501) begin
      mstatus <= _T_535;
    end else if (_T_429) begin
      mstatus <= _T_463;
    end
    if (reset) begin
      medeleg <= 64'h0;
    end else if (_T_393) begin
      medeleg <= _T_397;
    end
    if (reset) begin
      mideleg <= 64'h0;
    end else if (_T_561) begin
      mideleg <= _T_565;
    end
    if (reset) begin
      mscratch <= 64'h0;
    end else if (_T_579) begin
      mscratch <= wdata;
    end
    if (reset) begin
      pmpcfg0 <= 64'h0;
    end else if (_T_603) begin
      pmpcfg0 <= wdata;
    end
    if (reset) begin
      pmpcfg1 <= 64'h0;
    end else if (_T_573) begin
      pmpcfg1 <= wdata;
    end
    if (reset) begin
      pmpcfg2 <= 64'h0;
    end else if (_T_381) begin
      pmpcfg2 <= wdata;
    end
    if (reset) begin
      pmpcfg3 <= 64'h0;
    end else if (_T_555) begin
      pmpcfg3 <= wdata;
    end
    if (reset) begin
      pmpaddr0 <= 64'h0;
    end else if (_T_543) begin
      pmpaddr0 <= wdata;
    end
    if (reset) begin
      pmpaddr1 <= 64'h0;
    end else if (_T_375) begin
      pmpaddr1 <= wdata;
    end
    if (reset) begin
      pmpaddr2 <= 64'h0;
    end else if (_T_567) begin
      pmpaddr2 <= wdata;
    end
    if (reset) begin
      pmpaddr3 <= 64'h0;
    end else if (_T_483) begin
      pmpaddr3 <= wdata;
    end
    if (reset) begin
      stvec <= 64'h0;
    end else if (_T_399) begin
      stvec <= wdata;
    end
    if (reset) begin
      satp <= 64'h0;
    end else if (_T_369) begin
      satp <= wdata;
    end
    if (reset) begin
      sepc <= 64'h0;
    end else if (raiseExceptionIntr) begin
      if (delegS) begin
        sepc <= _T_772;
      end else if (_T_405) begin
        sepc <= wdata;
      end
    end else if (_T_405) begin
      sepc <= wdata;
    end
    if (reset) begin
      scause <= 64'h0;
    end else if (raiseExceptionIntr) begin
      if (delegS) begin
        scause <= causeNO;
      end else if (_T_609) begin
        scause <= wdata;
      end
    end else if (_T_609) begin
      scause <= wdata;
    end
    if (raiseExceptionIntr) begin
      if (delegS) begin
        if (tvalWen) begin
          stval <= 64'h0;
        end else if (_T_760) begin
          if (_T_779) begin
            if (_T_489) begin
              stval <= wdata;
            end
          end else if (hasInstrPageFault) begin
            if (io_cfIn_crossPageIPFFix) begin
              stval <= _T_767;
            end else begin
              stval <= _T_772;
            end
          end else begin
            stval <= _T_777;
          end
        end else if (_T_489) begin
          stval <= wdata;
        end
      end else if (_T_760) begin
        if (_T_779) begin
          if (_T_489) begin
            stval <= wdata;
          end
        end else begin
          stval <= _T_778;
        end
      end else if (_T_489) begin
        stval <= wdata;
      end
    end else if (_T_760) begin
      if (_T_779) begin
        stval <= _GEN_17;
      end else begin
        stval <= _T_778;
      end
    end else begin
      stval <= _GEN_17;
    end
    if (reset) begin
      sscratch <= 64'h0;
    end else if (_T_387) begin
      sscratch <= wdata;
    end
    if (reset) begin
      scounteren <= 64'h0;
    end else if (_T_597) begin
      scounteren <= wdata;
    end
    if (reset) begin
      lr <= 1'h0;
    end else if (_T_1308) begin
      lr <= 1'h0;
    end else if (_T_1229) begin
      lr <= 1'h0;
    end else if (set_lr) begin
      lr <= set_lr_val;
    end
    if (reset) begin
      lrAddr <= 64'h0;
    end else if (set_lr) begin
      lrAddr <= set_lr_addr;
    end
    if (reset) begin
      priviledgeMode <= 2'h3;
    end else if (raiseExceptionIntr) begin
      if (delegS) begin
        priviledgeMode <= 2'h1;
      end else begin
        priviledgeMode <= 2'h3;
      end
    end else if (_T_1388) begin
      priviledgeMode <= 2'h0;
    end else if (_T_1308) begin
      priviledgeMode <= _T_1363;
    end else if (_T_1229) begin
      priviledgeMode <= mstatusStruct_mpp;
    end
    if (reset) begin
      perfCnts_0 <= 64'h0;
    end else begin
      perfCnts_0 <= _T_1553;
    end
    if (reset) begin
      perfCnts_1 <= 64'h0;
    end else if (_T_477) begin
      perfCnts_1 <= wdata;
    end
    if (reset) begin
      perfCnts_2 <= 64'h0;
    end else if (perfCntCondMultiCommit) begin
      perfCnts_2 <= _T_1559;
    end else if (perfCntCondMinstret) begin
      perfCnts_2 <= _T_1557;
    end else if (_T_549) begin
      perfCnts_2 <= wdata;
    end
  end
endmodule
module MOU(
  input         io_in_valid,
  input  [6:0]  io_in_bits_func,
  input  [38:0] io_cfIn_pc,
  output [38:0] io_redirect_target,
  output        io_redirect_valid,
  output        flushICache_0,
  output        flushTLB_0
);
  wire  _T_2 = io_in_bits_func == 7'h1; // @[MOU.scala 52:36]
  wire  flushICache = io_in_valid & _T_2; // @[MOU.scala 52:27]
  wire  _T_12 = io_in_bits_func == 7'h2; // @[MOU.scala 56:33]
  wire  flushTLB = io_in_valid & _T_12; // @[MOU.scala 56:24]
  assign io_redirect_target = io_cfIn_pc + 39'h4; // @[MOU.scala 49:22]
  assign io_redirect_valid = io_in_valid; // @[MOU.scala 50:21]
  assign flushICache_0 = flushICache;
  assign flushTLB_0 = flushTLB;
endmodule
module EXU(
  input         clock,
  input         reset,
  output        io__in_ready,
  input         io__in_valid,
  input  [63:0] io__in_bits_cf_instr,
  input  [38:0] io__in_bits_cf_pc,
  input  [38:0] io__in_bits_cf_pnpc,
  input         io__in_bits_cf_exceptionVec_1,
  input         io__in_bits_cf_exceptionVec_2,
  input         io__in_bits_cf_exceptionVec_12,
  input         io__in_bits_cf_intrVec_0,
  input         io__in_bits_cf_intrVec_1,
  input         io__in_bits_cf_intrVec_2,
  input         io__in_bits_cf_intrVec_3,
  input         io__in_bits_cf_intrVec_4,
  input         io__in_bits_cf_intrVec_5,
  input         io__in_bits_cf_intrVec_6,
  input         io__in_bits_cf_intrVec_7,
  input         io__in_bits_cf_intrVec_8,
  input         io__in_bits_cf_intrVec_9,
  input         io__in_bits_cf_intrVec_10,
  input         io__in_bits_cf_intrVec_11,
  input  [3:0]  io__in_bits_cf_brIdx,
  input         io__in_bits_cf_crossPageIPFFix,
  input  [2:0]  io__in_bits_ctrl_fuType,
  input  [6:0]  io__in_bits_ctrl_fuOpType,
  input         io__in_bits_ctrl_rfWen,
  input  [4:0]  io__in_bits_ctrl_rfDest,
  input  [63:0] io__in_bits_data_src1,
  input  [63:0] io__in_bits_data_src2,
  input  [63:0] io__in_bits_data_imm,
  input         io__out_ready,
  output        io__out_valid,
  output [38:0] io__out_bits_decode_cf_pc,
  output [38:0] io__out_bits_decode_cf_redirect_target,
  output        io__out_bits_decode_cf_redirect_valid,
  output [2:0]  io__out_bits_decode_ctrl_fuType,
  output        io__out_bits_decode_ctrl_rfWen,
  output [4:0]  io__out_bits_decode_ctrl_rfDest,
  output [63:0] io__out_bits_commits_0,
  output [63:0] io__out_bits_commits_1,
  output [63:0] io__out_bits_commits_2,
  output [63:0] io__out_bits_commits_3,
  input         io__flush,
  input         io__dmem_req_ready,
  output        io__dmem_req_valid,
  output [38:0] io__dmem_req_bits_addr,
  output [2:0]  io__dmem_req_bits_size,
  output [3:0]  io__dmem_req_bits_cmd,
  output [7:0]  io__dmem_req_bits_wmask,
  output [63:0] io__dmem_req_bits_wdata,
  input         io__dmem_resp_valid,
  input  [63:0] io__dmem_resp_bits_rdata,
  output        io__forward_valid,
  output        io__forward_wb_rfWen,
  output [4:0]  io__forward_wb_rfDest,
  output [63:0] io__forward_wb_rfData,
  output [2:0]  io__forward_fuType,
  output [1:0]  io__memMMU_imem_priviledgeMode,
  output [1:0]  io__memMMU_dmem_priviledgeMode,
  output        io__memMMU_dmem_status_sum,
  output        io__memMMU_dmem_status_mxr,
  input         io__memMMU_dmem_loadPF,
  input         io__memMMU_dmem_storePF,
  input  [38:0] io__memMMU_dmem_addr,
  input         _T_38_0,
  output        flushICache,
  output [63:0] perfCnts_2,
  output [63:0] satp,
  output        _T_243_valid,
  output [38:0] _T_243_pc,
  output        _T_243_isMissPredict,
  output [38:0] _T_243_actualTarget,
  output        _T_243_actualTaken,
  output [6:0]  _T_243_fuOpType,
  output [1:0]  _T_243_btbType,
  output        _T_243_isRVC,
  input         io_in_valid,
  input         io_extra_mtip,
  output        amoReq,
  input         io_extra_meip_0,
  input         vmEnable,
  output [11:0] intrVec,
  input         _T_37_0,
  input         io_extra_msip,
  output        flushTLB,
  input         falseWire
);
  wire  alu_clock; // @[EXU.scala 45:19]
  wire  alu_reset; // @[EXU.scala 45:19]
  wire  alu_io_in_valid; // @[EXU.scala 45:19]
  wire [63:0] alu_io_in_bits_src1; // @[EXU.scala 45:19]
  wire [63:0] alu_io_in_bits_src2; // @[EXU.scala 45:19]
  wire [6:0] alu_io_in_bits_func; // @[EXU.scala 45:19]
  wire  alu_io_out_ready; // @[EXU.scala 45:19]
  wire  alu_io_out_valid; // @[EXU.scala 45:19]
  wire [63:0] alu_io_out_bits; // @[EXU.scala 45:19]
  wire [63:0] alu_io_cfIn_instr; // @[EXU.scala 45:19]
  wire [38:0] alu_io_cfIn_pc; // @[EXU.scala 45:19]
  wire [38:0] alu_io_cfIn_pnpc; // @[EXU.scala 45:19]
  wire [3:0] alu_io_cfIn_brIdx; // @[EXU.scala 45:19]
  wire [38:0] alu_io_redirect_target; // @[EXU.scala 45:19]
  wire  alu_io_redirect_valid; // @[EXU.scala 45:19]
  wire [63:0] alu_io_offset; // @[EXU.scala 45:19]
  wire  alu__T_243_0_valid; // @[EXU.scala 45:19]
  wire [38:0] alu__T_243_0_pc; // @[EXU.scala 45:19]
  wire  alu__T_243_0_isMissPredict; // @[EXU.scala 45:19]
  wire [38:0] alu__T_243_0_actualTarget; // @[EXU.scala 45:19]
  wire  alu__T_243_0_actualTaken; // @[EXU.scala 45:19]
  wire [6:0] alu__T_243_0_fuOpType; // @[EXU.scala 45:19]
  wire [1:0] alu__T_243_0_btbType; // @[EXU.scala 45:19]
  wire  alu__T_243_0_isRVC; // @[EXU.scala 45:19]
  wire  lsu_clock; // @[EXU.scala 53:19]
  wire  lsu_reset; // @[EXU.scala 53:19]
  wire  lsu_io__in_valid; // @[EXU.scala 53:19]
  wire [63:0] lsu_io__in_bits_src1; // @[EXU.scala 53:19]
  wire [63:0] lsu_io__in_bits_src2; // @[EXU.scala 53:19]
  wire [6:0] lsu_io__in_bits_func; // @[EXU.scala 53:19]
  wire  lsu_io__out_ready; // @[EXU.scala 53:19]
  wire  lsu_io__out_valid; // @[EXU.scala 53:19]
  wire [63:0] lsu_io__out_bits; // @[EXU.scala 53:19]
  wire [63:0] lsu_io__wdata; // @[EXU.scala 53:19]
  wire [31:0] lsu_io__instr; // @[EXU.scala 53:19]
  wire  lsu_io__dmem_req_ready; // @[EXU.scala 53:19]
  wire  lsu_io__dmem_req_valid; // @[EXU.scala 53:19]
  wire [38:0] lsu_io__dmem_req_bits_addr; // @[EXU.scala 53:19]
  wire [2:0] lsu_io__dmem_req_bits_size; // @[EXU.scala 53:19]
  wire [3:0] lsu_io__dmem_req_bits_cmd; // @[EXU.scala 53:19]
  wire [7:0] lsu_io__dmem_req_bits_wmask; // @[EXU.scala 53:19]
  wire [63:0] lsu_io__dmem_req_bits_wdata; // @[EXU.scala 53:19]
  wire  lsu_io__dmem_resp_valid; // @[EXU.scala 53:19]
  wire [63:0] lsu_io__dmem_resp_bits_rdata; // @[EXU.scala 53:19]
  wire  lsu_io__dtlbPF; // @[EXU.scala 53:19]
  wire  lsu_io__loadAddrMisaligned; // @[EXU.scala 53:19]
  wire  lsu_io__storeAddrMisaligned; // @[EXU.scala 53:19]
  wire  lsu_setLr_0; // @[EXU.scala 53:19]
  wire  lsu_DTLBPF; // @[EXU.scala 53:19]
  wire  lsu_amoReq_0; // @[EXU.scala 53:19]
  wire  lsu_DTLBENABLE; // @[EXU.scala 53:19]
  wire [63:0] lsu_io_in_bits_src1; // @[EXU.scala 53:19]
  wire  lsu_DTLBFINISH; // @[EXU.scala 53:19]
  wire [63:0] lsu_setLrAddr_0; // @[EXU.scala 53:19]
  wire  lsu_setLrVal_0; // @[EXU.scala 53:19]
  wire [63:0] lsu_lr_addr; // @[EXU.scala 53:19]
  wire  mdu_clock; // @[EXU.scala 62:19]
  wire  mdu_reset; // @[EXU.scala 62:19]
  wire  mdu_io_in_ready; // @[EXU.scala 62:19]
  wire  mdu_io_in_valid; // @[EXU.scala 62:19]
  wire [63:0] mdu_io_in_bits_src1; // @[EXU.scala 62:19]
  wire [63:0] mdu_io_in_bits_src2; // @[EXU.scala 62:19]
  wire [6:0] mdu_io_in_bits_func; // @[EXU.scala 62:19]
  wire  mdu_io_out_ready; // @[EXU.scala 62:19]
  wire  mdu_io_out_valid; // @[EXU.scala 62:19]
  wire [63:0] mdu_io_out_bits; // @[EXU.scala 62:19]
  wire  csr_clock; // @[EXU.scala 67:19]
  wire  csr_reset; // @[EXU.scala 67:19]
  wire  csr_io_in_valid; // @[EXU.scala 67:19]
  wire [63:0] csr_io_in_bits_src1; // @[EXU.scala 67:19]
  wire [63:0] csr_io_in_bits_src2; // @[EXU.scala 67:19]
  wire [6:0] csr_io_in_bits_func; // @[EXU.scala 67:19]
  wire  csr_io_out_ready; // @[EXU.scala 67:19]
  wire  csr_io_out_valid; // @[EXU.scala 67:19]
  wire [63:0] csr_io_out_bits; // @[EXU.scala 67:19]
  wire [63:0] csr_io_cfIn_instr; // @[EXU.scala 67:19]
  wire [38:0] csr_io_cfIn_pc; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_exceptionVec_1; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_exceptionVec_2; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_exceptionVec_4; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_exceptionVec_6; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_exceptionVec_12; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_intrVec_0; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_intrVec_1; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_intrVec_2; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_intrVec_3; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_intrVec_4; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_intrVec_5; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_intrVec_6; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_intrVec_7; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_intrVec_8; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_intrVec_9; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_intrVec_10; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_intrVec_11; // @[EXU.scala 67:19]
  wire  csr_io_cfIn_crossPageIPFFix; // @[EXU.scala 67:19]
  wire [38:0] csr_io_redirect_target; // @[EXU.scala 67:19]
  wire  csr_io_redirect_valid; // @[EXU.scala 67:19]
  wire  csr_io_instrValid; // @[EXU.scala 67:19]
  wire [1:0] csr_io_imemMMU_priviledgeMode; // @[EXU.scala 67:19]
  wire [1:0] csr_io_dmemMMU_priviledgeMode; // @[EXU.scala 67:19]
  wire  csr_io_dmemMMU_status_sum; // @[EXU.scala 67:19]
  wire  csr_io_dmemMMU_status_mxr; // @[EXU.scala 67:19]
  wire  csr_io_dmemMMU_loadPF; // @[EXU.scala 67:19]
  wire  csr_io_dmemMMU_storePF; // @[EXU.scala 67:19]
  wire [38:0] csr_io_dmemMMU_addr; // @[EXU.scala 67:19]
  wire  csr_io_wenFix; // @[EXU.scala 67:19]
  wire  csr_set_lr; // @[EXU.scala 67:19]
  wire [63:0] csr_perfCnts_2_0; // @[EXU.scala 67:19]
  wire [63:0] csr_satp_0; // @[EXU.scala 67:19]
  wire  csr_perfCntCondMinstret; // @[EXU.scala 67:19]
  wire  csr_mtip_0; // @[EXU.scala 67:19]
  wire  csr_meip_0; // @[EXU.scala 67:19]
  wire [63:0] csr_LSUADDR; // @[EXU.scala 67:19]
  wire [11:0] csr_intrVec_0; // @[EXU.scala 67:19]
  wire  csr_msip_0; // @[EXU.scala 67:19]
  wire [63:0] csr_set_lr_addr; // @[EXU.scala 67:19]
  wire  csr_perfCntCondMultiCommit; // @[EXU.scala 67:19]
  wire  csr_set_lr_val; // @[EXU.scala 67:19]
  wire [63:0] csr_lrAddr_0; // @[EXU.scala 67:19]
  wire  mou_io_in_valid; // @[EXU.scala 81:19]
  wire [6:0] mou_io_in_bits_func; // @[EXU.scala 81:19]
  wire [38:0] mou_io_cfIn_pc; // @[EXU.scala 81:19]
  wire [38:0] mou_io_redirect_target; // @[EXU.scala 81:19]
  wire  mou_io_redirect_valid; // @[EXU.scala 81:19]
  wire  mou_flushICache_0; // @[EXU.scala 81:19]
  wire  mou_flushTLB_0; // @[EXU.scala 81:19]
  wire  _T = io__in_bits_ctrl_fuType == 3'h0; // @[EXU.scala 43:57]
  wire  _T_1 = _T & io__in_valid; // @[EXU.scala 43:66]
  wire  _T_2 = ~io__flush; // @[EXU.scala 43:84]
  wire  _T_4 = io__in_bits_ctrl_fuType == 3'h1; // @[EXU.scala 43:57]
  wire  _T_5 = _T_4 & io__in_valid; // @[EXU.scala 43:66]
  wire  fuValids_1 = _T_5 & _T_2; // @[EXU.scala 43:81]
  wire  _T_8 = io__in_bits_ctrl_fuType == 3'h2; // @[EXU.scala 43:57]
  wire  _T_9 = _T_8 & io__in_valid; // @[EXU.scala 43:66]
  wire  _T_12 = io__in_bits_ctrl_fuType == 3'h3; // @[EXU.scala 43:57]
  wire  _T_13 = _T_12 & io__in_valid; // @[EXU.scala 43:66]
  wire  fuValids_3 = _T_13 & _T_2; // @[EXU.scala 43:81]
  wire  _T_16 = io__in_bits_ctrl_fuType == 3'h4; // @[EXU.scala 43:57]
  wire  _T_17 = _T_16 & io__in_valid; // @[EXU.scala 43:66]
  wire  lsuTlbPF = lsu_io__dtlbPF; // @[UnpipelinedLSU.scala 44:12]
  wire  _T_31 = ~lsuTlbPF; // @[EXU.scala 89:28]
  wire  _T_32 = ~lsu_io__loadAddrMisaligned; // @[EXU.scala 89:41]
  wire  _T_33 = _T_31 & _T_32; // @[EXU.scala 89:38]
  wire  _T_34 = ~lsu_io__storeAddrMisaligned; // @[EXU.scala 89:71]
  wire  _T_35 = _T_33 & _T_34; // @[EXU.scala 89:68]
  wire  _T_36 = ~fuValids_1; // @[EXU.scala 89:102]
  wire  _T_37 = _T_35 | _T_36; // @[EXU.scala 89:99]
  wire  _T_38 = io__in_bits_ctrl_rfWen & _T_37; // @[EXU.scala 89:24]
  wire  _T_39 = csr_io_wenFix & fuValids_3; // @[EXU.scala 89:144]
  wire  _T_40 = ~_T_39; // @[EXU.scala 89:128]
  wire [38:0] _T_42_target = csr_io_redirect_valid ? csr_io_redirect_target : alu_io_redirect_target; // @[EXU.scala 97:10]
  wire  _T_42_valid = csr_io_redirect_valid ? csr_io_redirect_valid : alu_io_redirect_valid; // @[EXU.scala 97:10]
  wire  _T_66 = 3'h1 == io__in_bits_ctrl_fuType; // @[Mux.scala 80:60]
  wire  _T_67 = _T_66 ? lsu_io__out_valid : 1'h1; // @[Mux.scala 80:57]
  wire  _T_68 = 3'h2 == io__in_bits_ctrl_fuType; // @[Mux.scala 80:60]
  wire  _T_69 = _T_68 ? mdu_io_out_valid : _T_67; // @[Mux.scala 80:57]
  wire  _T_71 = ~io__in_valid; // @[EXU.scala 114:18]
  wire  _T_74 = alu_io_out_ready & alu_io_out_valid; // @[Decoupled.scala 40:37]
  wire  isBru = io__in_bits_ctrl_fuOpType[4]; // @[ALU.scala 61:31]
  wire  _T_77 = ~isBru; // @[EXU.scala 123:46]
  wire  _T_78 = _T_74 & _T_77; // @[EXU.scala 123:43]
  wire  _T_80 = _T_74 & isBru; // @[EXU.scala 124:43]
  wire  _T_81 = lsu_io__out_ready & lsu_io__out_valid; // @[Decoupled.scala 40:37]
  wire  _T_82 = mdu_io_out_ready & mdu_io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_83 = csr_io_out_ready & csr_io_out_valid; // @[Decoupled.scala 40:37]
  ALU alu ( // @[EXU.scala 45:19]
    .clock(alu_clock),
    .reset(alu_reset),
    .io_in_valid(alu_io_in_valid),
    .io_in_bits_src1(alu_io_in_bits_src1),
    .io_in_bits_src2(alu_io_in_bits_src2),
    .io_in_bits_func(alu_io_in_bits_func),
    .io_out_ready(alu_io_out_ready),
    .io_out_valid(alu_io_out_valid),
    .io_out_bits(alu_io_out_bits),
    .io_cfIn_instr(alu_io_cfIn_instr),
    .io_cfIn_pc(alu_io_cfIn_pc),
    .io_cfIn_pnpc(alu_io_cfIn_pnpc),
    .io_cfIn_brIdx(alu_io_cfIn_brIdx),
    .io_redirect_target(alu_io_redirect_target),
    .io_redirect_valid(alu_io_redirect_valid),
    .io_offset(alu_io_offset),
    ._T_243_0_valid(alu__T_243_0_valid),
    ._T_243_0_pc(alu__T_243_0_pc),
    ._T_243_0_isMissPredict(alu__T_243_0_isMissPredict),
    ._T_243_0_actualTarget(alu__T_243_0_actualTarget),
    ._T_243_0_actualTaken(alu__T_243_0_actualTaken),
    ._T_243_0_fuOpType(alu__T_243_0_fuOpType),
    ._T_243_0_btbType(alu__T_243_0_btbType),
    ._T_243_0_isRVC(alu__T_243_0_isRVC)
  );
  UnpipelinedLSU lsu ( // @[EXU.scala 53:19]
    .clock(lsu_clock),
    .reset(lsu_reset),
    .io__in_valid(lsu_io__in_valid),
    .io__in_bits_src1(lsu_io__in_bits_src1),
    .io__in_bits_src2(lsu_io__in_bits_src2),
    .io__in_bits_func(lsu_io__in_bits_func),
    .io__out_ready(lsu_io__out_ready),
    .io__out_valid(lsu_io__out_valid),
    .io__out_bits(lsu_io__out_bits),
    .io__wdata(lsu_io__wdata),
    .io__instr(lsu_io__instr),
    .io__dmem_req_ready(lsu_io__dmem_req_ready),
    .io__dmem_req_valid(lsu_io__dmem_req_valid),
    .io__dmem_req_bits_addr(lsu_io__dmem_req_bits_addr),
    .io__dmem_req_bits_size(lsu_io__dmem_req_bits_size),
    .io__dmem_req_bits_cmd(lsu_io__dmem_req_bits_cmd),
    .io__dmem_req_bits_wmask(lsu_io__dmem_req_bits_wmask),
    .io__dmem_req_bits_wdata(lsu_io__dmem_req_bits_wdata),
    .io__dmem_resp_valid(lsu_io__dmem_resp_valid),
    .io__dmem_resp_bits_rdata(lsu_io__dmem_resp_bits_rdata),
    .io__dtlbPF(lsu_io__dtlbPF),
    .io__loadAddrMisaligned(lsu_io__loadAddrMisaligned),
    .io__storeAddrMisaligned(lsu_io__storeAddrMisaligned),
    .setLr_0(lsu_setLr_0),
    .DTLBPF(lsu_DTLBPF),
    .amoReq_0(lsu_amoReq_0),
    .DTLBENABLE(lsu_DTLBENABLE),
    .io_in_bits_src1(lsu_io_in_bits_src1),
    .DTLBFINISH(lsu_DTLBFINISH),
    .setLrAddr_0(lsu_setLrAddr_0),
    .setLrVal_0(lsu_setLrVal_0),
    .lr_addr(lsu_lr_addr)
  );
  MDU mdu ( // @[EXU.scala 62:19]
    .clock(mdu_clock),
    .reset(mdu_reset),
    .io_in_ready(mdu_io_in_ready),
    .io_in_valid(mdu_io_in_valid),
    .io_in_bits_src1(mdu_io_in_bits_src1),
    .io_in_bits_src2(mdu_io_in_bits_src2),
    .io_in_bits_func(mdu_io_in_bits_func),
    .io_out_ready(mdu_io_out_ready),
    .io_out_valid(mdu_io_out_valid),
    .io_out_bits(mdu_io_out_bits)
  );
  CSR csr ( // @[EXU.scala 67:19]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_in_valid(csr_io_in_valid),
    .io_in_bits_src1(csr_io_in_bits_src1),
    .io_in_bits_src2(csr_io_in_bits_src2),
    .io_in_bits_func(csr_io_in_bits_func),
    .io_out_ready(csr_io_out_ready),
    .io_out_valid(csr_io_out_valid),
    .io_out_bits(csr_io_out_bits),
    .io_cfIn_instr(csr_io_cfIn_instr),
    .io_cfIn_pc(csr_io_cfIn_pc),
    .io_cfIn_exceptionVec_1(csr_io_cfIn_exceptionVec_1),
    .io_cfIn_exceptionVec_2(csr_io_cfIn_exceptionVec_2),
    .io_cfIn_exceptionVec_4(csr_io_cfIn_exceptionVec_4),
    .io_cfIn_exceptionVec_6(csr_io_cfIn_exceptionVec_6),
    .io_cfIn_exceptionVec_12(csr_io_cfIn_exceptionVec_12),
    .io_cfIn_intrVec_0(csr_io_cfIn_intrVec_0),
    .io_cfIn_intrVec_1(csr_io_cfIn_intrVec_1),
    .io_cfIn_intrVec_2(csr_io_cfIn_intrVec_2),
    .io_cfIn_intrVec_3(csr_io_cfIn_intrVec_3),
    .io_cfIn_intrVec_4(csr_io_cfIn_intrVec_4),
    .io_cfIn_intrVec_5(csr_io_cfIn_intrVec_5),
    .io_cfIn_intrVec_6(csr_io_cfIn_intrVec_6),
    .io_cfIn_intrVec_7(csr_io_cfIn_intrVec_7),
    .io_cfIn_intrVec_8(csr_io_cfIn_intrVec_8),
    .io_cfIn_intrVec_9(csr_io_cfIn_intrVec_9),
    .io_cfIn_intrVec_10(csr_io_cfIn_intrVec_10),
    .io_cfIn_intrVec_11(csr_io_cfIn_intrVec_11),
    .io_cfIn_crossPageIPFFix(csr_io_cfIn_crossPageIPFFix),
    .io_redirect_target(csr_io_redirect_target),
    .io_redirect_valid(csr_io_redirect_valid),
    .io_instrValid(csr_io_instrValid),
    .io_imemMMU_priviledgeMode(csr_io_imemMMU_priviledgeMode),
    .io_dmemMMU_priviledgeMode(csr_io_dmemMMU_priviledgeMode),
    .io_dmemMMU_status_sum(csr_io_dmemMMU_status_sum),
    .io_dmemMMU_status_mxr(csr_io_dmemMMU_status_mxr),
    .io_dmemMMU_loadPF(csr_io_dmemMMU_loadPF),
    .io_dmemMMU_storePF(csr_io_dmemMMU_storePF),
    .io_dmemMMU_addr(csr_io_dmemMMU_addr),
    .io_wenFix(csr_io_wenFix),
    .set_lr(csr_set_lr),
    .perfCnts_2_0(csr_perfCnts_2_0),
    .satp_0(csr_satp_0),
    .perfCntCondMinstret(csr_perfCntCondMinstret),
    .mtip_0(csr_mtip_0),
    .meip_0(csr_meip_0),
    .LSUADDR(csr_LSUADDR),
    .intrVec_0(csr_intrVec_0),
    .msip_0(csr_msip_0),
    .set_lr_addr(csr_set_lr_addr),
    .perfCntCondMultiCommit(csr_perfCntCondMultiCommit),
    .set_lr_val(csr_set_lr_val),
    .lrAddr_0(csr_lrAddr_0)
  );
  MOU mou ( // @[EXU.scala 81:19]
    .io_in_valid(mou_io_in_valid),
    .io_in_bits_func(mou_io_in_bits_func),
    .io_cfIn_pc(mou_io_cfIn_pc),
    .io_redirect_target(mou_io_redirect_target),
    .io_redirect_valid(mou_io_redirect_valid),
    .flushICache_0(mou_flushICache_0),
    .flushTLB_0(mou_flushTLB_0)
  );
  assign io__in_ready = _T_71 | io__out_valid; // @[EXU.scala 114:15]
  assign io__out_valid = io__in_valid & _T_69; // @[EXU.scala 103:16]
  assign io__out_bits_decode_cf_pc = io__in_bits_cf_pc; // @[EXU.scala 93:28]
  assign io__out_bits_decode_cf_redirect_target = mou_io_redirect_valid ? mou_io_redirect_target : _T_42_target; // @[EXU.scala 95:34]
  assign io__out_bits_decode_cf_redirect_valid = mou_io_redirect_valid ? mou_io_redirect_valid : _T_42_valid; // @[EXU.scala 95:34]
  assign io__out_bits_decode_ctrl_fuType = io__in_bits_ctrl_fuType; // @[EXU.scala 91:14]
  assign io__out_bits_decode_ctrl_rfWen = _T_38 & _T_40; // @[EXU.scala 89:13]
  assign io__out_bits_decode_ctrl_rfDest = io__in_bits_ctrl_rfDest; // @[EXU.scala 90:14]
  assign io__out_bits_commits_0 = alu_io_out_bits; // @[EXU.scala 108:35]
  assign io__out_bits_commits_1 = lsu_io__out_bits; // @[EXU.scala 109:35]
  assign io__out_bits_commits_2 = mdu_io_out_bits; // @[EXU.scala 111:35]
  assign io__out_bits_commits_3 = csr_io_out_bits; // @[EXU.scala 110:35]
  assign io__dmem_req_valid = lsu_io__dmem_req_valid; // @[EXU.scala 59:11]
  assign io__dmem_req_bits_addr = lsu_io__dmem_req_bits_addr; // @[EXU.scala 59:11]
  assign io__dmem_req_bits_size = lsu_io__dmem_req_bits_size; // @[EXU.scala 59:11]
  assign io__dmem_req_bits_cmd = lsu_io__dmem_req_bits_cmd; // @[EXU.scala 59:11]
  assign io__dmem_req_bits_wmask = lsu_io__dmem_req_bits_wmask; // @[EXU.scala 59:11]
  assign io__dmem_req_bits_wdata = lsu_io__dmem_req_bits_wdata; // @[EXU.scala 59:11]
  assign io__forward_valid = io__in_valid; // @[EXU.scala 116:20]
  assign io__forward_wb_rfWen = io__in_bits_ctrl_rfWen; // @[EXU.scala 117:23]
  assign io__forward_wb_rfDest = io__in_bits_ctrl_rfDest; // @[EXU.scala 118:24]
  assign io__forward_wb_rfData = _T_74 ? alu_io_out_bits : lsu_io__out_bits; // @[EXU.scala 119:24]
  assign io__forward_fuType = io__in_bits_ctrl_fuType; // @[EXU.scala 120:21]
  assign io__memMMU_imem_priviledgeMode = csr_io_imemMMU_priviledgeMode; // @[EXU.scala 78:18]
  assign io__memMMU_dmem_priviledgeMode = csr_io_dmemMMU_priviledgeMode; // @[EXU.scala 79:18]
  assign io__memMMU_dmem_status_sum = csr_io_dmemMMU_status_sum; // @[EXU.scala 79:18]
  assign io__memMMU_dmem_status_mxr = csr_io_dmemMMU_status_mxr; // @[EXU.scala 79:18]
  assign flushICache = mou_flushICache_0;
  assign perfCnts_2 = csr_perfCnts_2_0;
  assign satp = csr_satp_0;
  assign _T_243_valid = alu__T_243_0_valid;
  assign _T_243_pc = alu__T_243_0_pc;
  assign _T_243_isMissPredict = alu__T_243_0_isMissPredict;
  assign _T_243_actualTarget = alu__T_243_0_actualTarget;
  assign _T_243_actualTaken = alu__T_243_0_actualTaken;
  assign _T_243_fuOpType = alu__T_243_0_fuOpType;
  assign _T_243_btbType = alu__T_243_0_btbType;
  assign _T_243_isRVC = alu__T_243_0_isRVC;
  assign amoReq = lsu_amoReq_0;
  assign intrVec = csr_intrVec_0;
  assign flushTLB = mou_flushTLB_0;
  assign alu_clock = clock;
  assign alu_reset = reset;
  assign alu_io_in_valid = _T_1 & _T_2; // @[ALU.scala 79:16]
  assign alu_io_in_bits_src1 = io__in_bits_data_src1; // @[ALU.scala 80:15]
  assign alu_io_in_bits_src2 = io__in_bits_data_src2; // @[ALU.scala 81:15]
  assign alu_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[ALU.scala 82:15]
  assign alu_io_out_ready = 1'h1; // @[EXU.scala 49:20]
  assign alu_io_cfIn_instr = io__in_bits_cf_instr; // @[EXU.scala 47:15]
  assign alu_io_cfIn_pc = io__in_bits_cf_pc; // @[EXU.scala 47:15]
  assign alu_io_cfIn_pnpc = io__in_bits_cf_pnpc; // @[EXU.scala 47:15]
  assign alu_io_cfIn_brIdx = io__in_bits_cf_brIdx; // @[EXU.scala 47:15]
  assign alu_io_offset = io__in_bits_data_imm; // @[EXU.scala 48:17]
  assign lsu_clock = clock;
  assign lsu_reset = reset;
  assign lsu_io__in_valid = _T_5 & _T_2; // @[UnpipelinedLSU.scala 40:16]
  assign lsu_io__in_bits_src1 = io__in_bits_data_src1; // @[UnpipelinedLSU.scala 41:15]
  assign lsu_io__in_bits_src2 = io__in_bits_data_imm; // @[UnpipelinedLSU.scala 42:15]
  assign lsu_io__in_bits_func = io__in_bits_ctrl_fuOpType; // @[UnpipelinedLSU.scala 43:15]
  assign lsu_io__out_ready = 1'h1; // @[EXU.scala 60:20]
  assign lsu_io__wdata = io__in_bits_data_src2; // @[EXU.scala 56:16]
  assign lsu_io__instr = io__in_bits_cf_instr[31:0]; // @[EXU.scala 57:16]
  assign lsu_io__dmem_req_ready = io__dmem_req_ready; // @[EXU.scala 59:11]
  assign lsu_io__dmem_resp_valid = io__dmem_resp_valid; // @[EXU.scala 59:11]
  assign lsu_io__dmem_resp_bits_rdata = io__dmem_resp_bits_rdata; // @[EXU.scala 59:11]
  assign lsu_DTLBPF = _T_38_0;
  assign lsu_DTLBENABLE = vmEnable;
  assign lsu_DTLBFINISH = _T_37_0;
  assign lsu_lr_addr = csr_lrAddr_0;
  assign mdu_clock = clock;
  assign mdu_reset = reset;
  assign mdu_io_in_valid = _T_9 & _T_2; // @[MDU.scala 140:16]
  assign mdu_io_in_bits_src1 = io__in_bits_data_src1; // @[MDU.scala 141:15]
  assign mdu_io_in_bits_src2 = io__in_bits_data_src2; // @[MDU.scala 142:15]
  assign mdu_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[MDU.scala 143:15]
  assign mdu_io_out_ready = 1'h1; // @[EXU.scala 64:20]
  assign csr_clock = clock;
  assign csr_reset = reset;
  assign csr_io_in_valid = _T_13 & _T_2; // @[CSR.scala 196:16]
  assign csr_io_in_bits_src1 = io__in_bits_data_src1; // @[CSR.scala 197:15]
  assign csr_io_in_bits_src2 = io__in_bits_data_src2; // @[CSR.scala 198:15]
  assign csr_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[CSR.scala 199:15]
  assign csr_io_out_ready = 1'h1; // @[EXU.scala 76:20]
  assign csr_io_cfIn_instr = io__in_bits_cf_instr; // @[EXU.scala 69:15]
  assign csr_io_cfIn_pc = io__in_bits_cf_pc; // @[EXU.scala 69:15]
  assign csr_io_cfIn_exceptionVec_1 = io__in_bits_cf_exceptionVec_1; // @[EXU.scala 69:15]
  assign csr_io_cfIn_exceptionVec_2 = io__in_bits_cf_exceptionVec_2; // @[EXU.scala 69:15]
  assign csr_io_cfIn_exceptionVec_4 = lsu_io__loadAddrMisaligned; // @[EXU.scala 69:15 EXU.scala 70:48]
  assign csr_io_cfIn_exceptionVec_6 = lsu_io__storeAddrMisaligned; // @[EXU.scala 69:15 EXU.scala 71:49]
  assign csr_io_cfIn_exceptionVec_12 = io__in_bits_cf_exceptionVec_12; // @[EXU.scala 69:15]
  assign csr_io_cfIn_intrVec_0 = io__in_bits_cf_intrVec_0; // @[EXU.scala 69:15]
  assign csr_io_cfIn_intrVec_1 = io__in_bits_cf_intrVec_1; // @[EXU.scala 69:15]
  assign csr_io_cfIn_intrVec_2 = io__in_bits_cf_intrVec_2; // @[EXU.scala 69:15]
  assign csr_io_cfIn_intrVec_3 = io__in_bits_cf_intrVec_3; // @[EXU.scala 69:15]
  assign csr_io_cfIn_intrVec_4 = io__in_bits_cf_intrVec_4; // @[EXU.scala 69:15]
  assign csr_io_cfIn_intrVec_5 = io__in_bits_cf_intrVec_5; // @[EXU.scala 69:15]
  assign csr_io_cfIn_intrVec_6 = io__in_bits_cf_intrVec_6; // @[EXU.scala 69:15]
  assign csr_io_cfIn_intrVec_7 = io__in_bits_cf_intrVec_7; // @[EXU.scala 69:15]
  assign csr_io_cfIn_intrVec_8 = io__in_bits_cf_intrVec_8; // @[EXU.scala 69:15]
  assign csr_io_cfIn_intrVec_9 = io__in_bits_cf_intrVec_9; // @[EXU.scala 69:15]
  assign csr_io_cfIn_intrVec_10 = io__in_bits_cf_intrVec_10; // @[EXU.scala 69:15]
  assign csr_io_cfIn_intrVec_11 = io__in_bits_cf_intrVec_11; // @[EXU.scala 69:15]
  assign csr_io_cfIn_crossPageIPFFix = io__in_bits_cf_crossPageIPFFix; // @[EXU.scala 69:15]
  assign csr_io_instrValid = io__in_valid & _T_2; // @[EXU.scala 72:21]
  assign csr_io_dmemMMU_loadPF = io__memMMU_dmem_loadPF; // @[EXU.scala 79:18]
  assign csr_io_dmemMMU_storePF = io__memMMU_dmem_storePF; // @[EXU.scala 79:18]
  assign csr_io_dmemMMU_addr = io__memMMU_dmem_addr; // @[EXU.scala 79:18]
  assign csr_set_lr = lsu_setLr_0;
  assign csr_perfCntCondMinstret = io_in_valid;
  assign csr_mtip_0 = io_extra_mtip;
  assign csr_meip_0 = io_extra_meip_0;
  assign csr_LSUADDR = lsu_io_in_bits_src1;
  assign csr_msip_0 = io_extra_msip;
  assign csr_set_lr_addr = lsu_setLrAddr_0;
  assign csr_perfCntCondMultiCommit = falseWire;
  assign csr_set_lr_val = lsu_setLrVal_0;
  assign mou_io_in_valid = _T_17 & _T_2; // @[MOU.scala 42:16]
  assign mou_io_in_bits_func = io__in_bits_ctrl_fuOpType; // @[MOU.scala 45:15]
  assign mou_io_cfIn_pc = io__in_bits_cf_pc; // @[EXU.scala 84:15]
endmodule
module WBU(
  input         io__in_valid,
  input  [38:0] io__in_bits_decode_cf_pc,
  input  [38:0] io__in_bits_decode_cf_redirect_target,
  input         io__in_bits_decode_cf_redirect_valid,
  input  [2:0]  io__in_bits_decode_ctrl_fuType,
  input         io__in_bits_decode_ctrl_rfWen,
  input  [4:0]  io__in_bits_decode_ctrl_rfDest,
  input  [63:0] io__in_bits_commits_0,
  input  [63:0] io__in_bits_commits_1,
  input  [63:0] io__in_bits_commits_2,
  input  [63:0] io__in_bits_commits_3,
  output        io__wb_rfWen,
  output [4:0]  io__wb_rfDest,
  output [63:0] io__wb_rfData,
  output [38:0] io__redirect_target,
  output        io__redirect_valid,
  output [38:0] io_in_bits_decode_cf_pc,
  output [4:0]  io_wb_rfDest,
  output        io_in_valid,
  output        io_wb_rfWen,
  output [63:0] io_wb_rfData,
  output        io_in_valid_0,
  output        falseWire_0
);
  wire [63:0] _GEN_1 = 3'h1 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_1 : io__in_bits_commits_0; // @[WBU.scala 33:16]
  wire [63:0] _GEN_2 = 3'h2 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_2 : _GEN_1; // @[WBU.scala 33:16]
  wire [63:0] _GEN_3 = 3'h3 == io__in_bits_decode_ctrl_fuType ? io__in_bits_commits_3 : _GEN_2; // @[WBU.scala 33:16]
  wire  _T_5 = 1'h0;
  wire  falseWire = 1'h0;
  assign io__wb_rfWen = io__in_bits_decode_ctrl_rfWen & io__in_valid; // @[WBU.scala 31:15]
  assign io__wb_rfDest = io__in_bits_decode_ctrl_rfDest; // @[WBU.scala 32:16]
  assign io__wb_rfData = 3'h4 == io__in_bits_decode_ctrl_fuType ? 64'h0 : _GEN_3; // @[WBU.scala 33:16]
  assign io__redirect_target = io__in_bits_decode_cf_redirect_target; // @[WBU.scala 37:15]
  assign io__redirect_valid = io__in_bits_decode_cf_redirect_valid & io__in_valid; // @[WBU.scala 37:15 WBU.scala 38:21]
  assign io_in_bits_decode_cf_pc = io__in_bits_decode_cf_pc;
  assign io_wb_rfDest = io__wb_rfDest;
  assign io_in_valid = io__in_valid;
  assign io_wb_rfWen = io__wb_rfWen;
  assign io_wb_rfData = io__wb_rfData;
  assign io_in_valid_0 = io__in_valid;
  assign falseWire_0 = _T_5;
endmodule
module Backend_inorder(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [63:0] io_in_0_bits_cf_instr,
  input  [38:0] io_in_0_bits_cf_pc,
  input  [38:0] io_in_0_bits_cf_pnpc,
  input         io_in_0_bits_cf_exceptionVec_1,
  input         io_in_0_bits_cf_exceptionVec_2,
  input         io_in_0_bits_cf_exceptionVec_12,
  input         io_in_0_bits_cf_intrVec_0,
  input         io_in_0_bits_cf_intrVec_1,
  input         io_in_0_bits_cf_intrVec_2,
  input         io_in_0_bits_cf_intrVec_3,
  input         io_in_0_bits_cf_intrVec_4,
  input         io_in_0_bits_cf_intrVec_5,
  input         io_in_0_bits_cf_intrVec_6,
  input         io_in_0_bits_cf_intrVec_7,
  input         io_in_0_bits_cf_intrVec_8,
  input         io_in_0_bits_cf_intrVec_9,
  input         io_in_0_bits_cf_intrVec_10,
  input         io_in_0_bits_cf_intrVec_11,
  input  [3:0]  io_in_0_bits_cf_brIdx,
  input         io_in_0_bits_cf_crossPageIPFFix,
  input         io_in_0_bits_ctrl_src1Type,
  input         io_in_0_bits_ctrl_src2Type,
  input  [2:0]  io_in_0_bits_ctrl_fuType,
  input  [6:0]  io_in_0_bits_ctrl_fuOpType,
  input  [4:0]  io_in_0_bits_ctrl_rfSrc1,
  input  [4:0]  io_in_0_bits_ctrl_rfSrc2,
  input         io_in_0_bits_ctrl_rfWen,
  input  [4:0]  io_in_0_bits_ctrl_rfDest,
  input  [63:0] io_in_0_bits_data_imm,
  input  [1:0]  io_flush,
  input         io_dmem_req_ready,
  output        io_dmem_req_valid,
  output [38:0] io_dmem_req_bits_addr,
  output [2:0]  io_dmem_req_bits_size,
  output [3:0]  io_dmem_req_bits_cmd,
  output [7:0]  io_dmem_req_bits_wmask,
  output [63:0] io_dmem_req_bits_wdata,
  input         io_dmem_resp_valid,
  input  [63:0] io_dmem_resp_bits_rdata,
  output [1:0]  io_memMMU_imem_priviledgeMode,
  output [1:0]  io_memMMU_dmem_priviledgeMode,
  output        io_memMMU_dmem_status_sum,
  output        io_memMMU_dmem_status_mxr,
  input         io_memMMU_dmem_loadPF,
  input         io_memMMU_dmem_storePF,
  input  [38:0] io_memMMU_dmem_addr,
  output [38:0] io_redirect_target,
  output        io_redirect_valid,
  input         _T_38,
  output        flushICache,
  output [63:0] perfCnts_2,
  output [38:0] io_in_bits_decode_cf_pc,
  output [63:0] satp,
  output        _T_243_valid,
  output [38:0] _T_243_pc,
  output        _T_243_isMissPredict,
  output [38:0] _T_243_actualTarget,
  output        _T_243_actualTaken,
  output [6:0]  _T_243_fuOpType,
  output [1:0]  _T_243_btbType,
  output        _T_243_isRVC,
  output [4:0]  io_wb_rfDest,
  input         io_extra_mtip,
  output        amoReq,
  input         io_extra_meip_0,
  input         vmEnable,
  output        io_wb_rfWen,
  output [63:0] io_wb_rfData,
  output [11:0] intrVec,
  input         _T_37,
  input         io_extra_msip,
  output        flushTLB,
  output        io_in_valid_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [63:0] _RAND_35;
  reg [63:0] _RAND_36;
  reg [63:0] _RAND_37;
  reg [63:0] _RAND_38;
`endif // RANDOMIZE_REG_INIT
  wire  isu_clock; // @[Backend.scala 675:20]
  wire  isu_reset; // @[Backend.scala 675:20]
  wire  isu_io_in_0_ready; // @[Backend.scala 675:20]
  wire  isu_io_in_0_valid; // @[Backend.scala 675:20]
  wire [63:0] isu_io_in_0_bits_cf_instr; // @[Backend.scala 675:20]
  wire [38:0] isu_io_in_0_bits_cf_pc; // @[Backend.scala 675:20]
  wire [38:0] isu_io_in_0_bits_cf_pnpc; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_1; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_2; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_exceptionVec_12; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_intrVec_0; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_intrVec_1; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_intrVec_2; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_intrVec_3; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_intrVec_4; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_intrVec_5; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_intrVec_6; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_intrVec_7; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_intrVec_8; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_intrVec_9; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_intrVec_10; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_intrVec_11; // @[Backend.scala 675:20]
  wire [3:0] isu_io_in_0_bits_cf_brIdx; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_cf_crossPageIPFFix; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_ctrl_src1Type; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_ctrl_src2Type; // @[Backend.scala 675:20]
  wire [2:0] isu_io_in_0_bits_ctrl_fuType; // @[Backend.scala 675:20]
  wire [6:0] isu_io_in_0_bits_ctrl_fuOpType; // @[Backend.scala 675:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfSrc1; // @[Backend.scala 675:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfSrc2; // @[Backend.scala 675:20]
  wire  isu_io_in_0_bits_ctrl_rfWen; // @[Backend.scala 675:20]
  wire [4:0] isu_io_in_0_bits_ctrl_rfDest; // @[Backend.scala 675:20]
  wire [63:0] isu_io_in_0_bits_data_imm; // @[Backend.scala 675:20]
  wire  isu_io_out_ready; // @[Backend.scala 675:20]
  wire  isu_io_out_valid; // @[Backend.scala 675:20]
  wire [63:0] isu_io_out_bits_cf_instr; // @[Backend.scala 675:20]
  wire [38:0] isu_io_out_bits_cf_pc; // @[Backend.scala 675:20]
  wire [38:0] isu_io_out_bits_cf_pnpc; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_exceptionVec_1; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_exceptionVec_2; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_exceptionVec_12; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_intrVec_0; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_intrVec_1; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_intrVec_2; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_intrVec_3; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_intrVec_4; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_intrVec_5; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_intrVec_6; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_intrVec_7; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_intrVec_8; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_intrVec_9; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_intrVec_10; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_intrVec_11; // @[Backend.scala 675:20]
  wire [3:0] isu_io_out_bits_cf_brIdx; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_cf_crossPageIPFFix; // @[Backend.scala 675:20]
  wire [2:0] isu_io_out_bits_ctrl_fuType; // @[Backend.scala 675:20]
  wire [6:0] isu_io_out_bits_ctrl_fuOpType; // @[Backend.scala 675:20]
  wire  isu_io_out_bits_ctrl_rfWen; // @[Backend.scala 675:20]
  wire [4:0] isu_io_out_bits_ctrl_rfDest; // @[Backend.scala 675:20]
  wire [63:0] isu_io_out_bits_data_src1; // @[Backend.scala 675:20]
  wire [63:0] isu_io_out_bits_data_src2; // @[Backend.scala 675:20]
  wire [63:0] isu_io_out_bits_data_imm; // @[Backend.scala 675:20]
  wire  isu_io_wb_rfWen; // @[Backend.scala 675:20]
  wire [4:0] isu_io_wb_rfDest; // @[Backend.scala 675:20]
  wire [63:0] isu_io_wb_rfData; // @[Backend.scala 675:20]
  wire  isu_io_forward_valid; // @[Backend.scala 675:20]
  wire  isu_io_forward_wb_rfWen; // @[Backend.scala 675:20]
  wire [4:0] isu_io_forward_wb_rfDest; // @[Backend.scala 675:20]
  wire [63:0] isu_io_forward_wb_rfData; // @[Backend.scala 675:20]
  wire [2:0] isu_io_forward_fuType; // @[Backend.scala 675:20]
  wire  isu_io_flush; // @[Backend.scala 675:20]
  wire  exu_clock; // @[Backend.scala 676:20]
  wire  exu_reset; // @[Backend.scala 676:20]
  wire  exu_io__in_ready; // @[Backend.scala 676:20]
  wire  exu_io__in_valid; // @[Backend.scala 676:20]
  wire [63:0] exu_io__in_bits_cf_instr; // @[Backend.scala 676:20]
  wire [38:0] exu_io__in_bits_cf_pc; // @[Backend.scala 676:20]
  wire [38:0] exu_io__in_bits_cf_pnpc; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_exceptionVec_1; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_exceptionVec_2; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_exceptionVec_12; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_intrVec_0; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_intrVec_1; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_intrVec_2; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_intrVec_3; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_intrVec_4; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_intrVec_5; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_intrVec_6; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_intrVec_7; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_intrVec_8; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_intrVec_9; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_intrVec_10; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_intrVec_11; // @[Backend.scala 676:20]
  wire [3:0] exu_io__in_bits_cf_brIdx; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_cf_crossPageIPFFix; // @[Backend.scala 676:20]
  wire [2:0] exu_io__in_bits_ctrl_fuType; // @[Backend.scala 676:20]
  wire [6:0] exu_io__in_bits_ctrl_fuOpType; // @[Backend.scala 676:20]
  wire  exu_io__in_bits_ctrl_rfWen; // @[Backend.scala 676:20]
  wire [4:0] exu_io__in_bits_ctrl_rfDest; // @[Backend.scala 676:20]
  wire [63:0] exu_io__in_bits_data_src1; // @[Backend.scala 676:20]
  wire [63:0] exu_io__in_bits_data_src2; // @[Backend.scala 676:20]
  wire [63:0] exu_io__in_bits_data_imm; // @[Backend.scala 676:20]
  wire  exu_io__out_ready; // @[Backend.scala 676:20]
  wire  exu_io__out_valid; // @[Backend.scala 676:20]
  wire [38:0] exu_io__out_bits_decode_cf_pc; // @[Backend.scala 676:20]
  wire [38:0] exu_io__out_bits_decode_cf_redirect_target; // @[Backend.scala 676:20]
  wire  exu_io__out_bits_decode_cf_redirect_valid; // @[Backend.scala 676:20]
  wire [2:0] exu_io__out_bits_decode_ctrl_fuType; // @[Backend.scala 676:20]
  wire  exu_io__out_bits_decode_ctrl_rfWen; // @[Backend.scala 676:20]
  wire [4:0] exu_io__out_bits_decode_ctrl_rfDest; // @[Backend.scala 676:20]
  wire [63:0] exu_io__out_bits_commits_0; // @[Backend.scala 676:20]
  wire [63:0] exu_io__out_bits_commits_1; // @[Backend.scala 676:20]
  wire [63:0] exu_io__out_bits_commits_2; // @[Backend.scala 676:20]
  wire [63:0] exu_io__out_bits_commits_3; // @[Backend.scala 676:20]
  wire  exu_io__flush; // @[Backend.scala 676:20]
  wire  exu_io__dmem_req_ready; // @[Backend.scala 676:20]
  wire  exu_io__dmem_req_valid; // @[Backend.scala 676:20]
  wire [38:0] exu_io__dmem_req_bits_addr; // @[Backend.scala 676:20]
  wire [2:0] exu_io__dmem_req_bits_size; // @[Backend.scala 676:20]
  wire [3:0] exu_io__dmem_req_bits_cmd; // @[Backend.scala 676:20]
  wire [7:0] exu_io__dmem_req_bits_wmask; // @[Backend.scala 676:20]
  wire [63:0] exu_io__dmem_req_bits_wdata; // @[Backend.scala 676:20]
  wire  exu_io__dmem_resp_valid; // @[Backend.scala 676:20]
  wire [63:0] exu_io__dmem_resp_bits_rdata; // @[Backend.scala 676:20]
  wire  exu_io__forward_valid; // @[Backend.scala 676:20]
  wire  exu_io__forward_wb_rfWen; // @[Backend.scala 676:20]
  wire [4:0] exu_io__forward_wb_rfDest; // @[Backend.scala 676:20]
  wire [63:0] exu_io__forward_wb_rfData; // @[Backend.scala 676:20]
  wire [2:0] exu_io__forward_fuType; // @[Backend.scala 676:20]
  wire [1:0] exu_io__memMMU_imem_priviledgeMode; // @[Backend.scala 676:20]
  wire [1:0] exu_io__memMMU_dmem_priviledgeMode; // @[Backend.scala 676:20]
  wire  exu_io__memMMU_dmem_status_sum; // @[Backend.scala 676:20]
  wire  exu_io__memMMU_dmem_status_mxr; // @[Backend.scala 676:20]
  wire  exu_io__memMMU_dmem_loadPF; // @[Backend.scala 676:20]
  wire  exu_io__memMMU_dmem_storePF; // @[Backend.scala 676:20]
  wire [38:0] exu_io__memMMU_dmem_addr; // @[Backend.scala 676:20]
  wire  exu__T_38_0; // @[Backend.scala 676:20]
  wire  exu_flushICache; // @[Backend.scala 676:20]
  wire [63:0] exu_perfCnts_2; // @[Backend.scala 676:20]
  wire [63:0] exu_satp; // @[Backend.scala 676:20]
  wire  exu__T_243_valid; // @[Backend.scala 676:20]
  wire [38:0] exu__T_243_pc; // @[Backend.scala 676:20]
  wire  exu__T_243_isMissPredict; // @[Backend.scala 676:20]
  wire [38:0] exu__T_243_actualTarget; // @[Backend.scala 676:20]
  wire  exu__T_243_actualTaken; // @[Backend.scala 676:20]
  wire [6:0] exu__T_243_fuOpType; // @[Backend.scala 676:20]
  wire [1:0] exu__T_243_btbType; // @[Backend.scala 676:20]
  wire  exu__T_243_isRVC; // @[Backend.scala 676:20]
  wire  exu_io_in_valid; // @[Backend.scala 676:20]
  wire  exu_io_extra_mtip; // @[Backend.scala 676:20]
  wire  exu_amoReq; // @[Backend.scala 676:20]
  wire  exu_io_extra_meip_0; // @[Backend.scala 676:20]
  wire  exu_vmEnable; // @[Backend.scala 676:20]
  wire [11:0] exu_intrVec; // @[Backend.scala 676:20]
  wire  exu__T_37_0; // @[Backend.scala 676:20]
  wire  exu_io_extra_msip; // @[Backend.scala 676:20]
  wire  exu_flushTLB; // @[Backend.scala 676:20]
  wire  exu_falseWire; // @[Backend.scala 676:20]
  wire  wbu_io__in_valid; // @[Backend.scala 677:20]
  wire [38:0] wbu_io__in_bits_decode_cf_pc; // @[Backend.scala 677:20]
  wire [38:0] wbu_io__in_bits_decode_cf_redirect_target; // @[Backend.scala 677:20]
  wire  wbu_io__in_bits_decode_cf_redirect_valid; // @[Backend.scala 677:20]
  wire [2:0] wbu_io__in_bits_decode_ctrl_fuType; // @[Backend.scala 677:20]
  wire  wbu_io__in_bits_decode_ctrl_rfWen; // @[Backend.scala 677:20]
  wire [4:0] wbu_io__in_bits_decode_ctrl_rfDest; // @[Backend.scala 677:20]
  wire [63:0] wbu_io__in_bits_commits_0; // @[Backend.scala 677:20]
  wire [63:0] wbu_io__in_bits_commits_1; // @[Backend.scala 677:20]
  wire [63:0] wbu_io__in_bits_commits_2; // @[Backend.scala 677:20]
  wire [63:0] wbu_io__in_bits_commits_3; // @[Backend.scala 677:20]
  wire  wbu_io__wb_rfWen; // @[Backend.scala 677:20]
  wire [4:0] wbu_io__wb_rfDest; // @[Backend.scala 677:20]
  wire [63:0] wbu_io__wb_rfData; // @[Backend.scala 677:20]
  wire [38:0] wbu_io__redirect_target; // @[Backend.scala 677:20]
  wire  wbu_io__redirect_valid; // @[Backend.scala 677:20]
  wire [38:0] wbu_io_in_bits_decode_cf_pc; // @[Backend.scala 677:20]
  wire [4:0] wbu_io_wb_rfDest; // @[Backend.scala 677:20]
  wire  wbu_io_in_valid; // @[Backend.scala 677:20]
  wire  wbu_io_wb_rfWen; // @[Backend.scala 677:20]
  wire [63:0] wbu_io_wb_rfData; // @[Backend.scala 677:20]
  wire  wbu_io_in_valid_0; // @[Backend.scala 677:20]
  wire  wbu_falseWire_0; // @[Backend.scala 677:20]
  wire  _T = exu_io__out_ready & exu_io__out_valid; // @[Decoupled.scala 40:37]
  reg  _T_2; // @[Pipeline.scala 24:24]
  wire  _GEN_0 = _T ? 1'h0 : _T_2; // @[Pipeline.scala 25:25]
  wire  _T_3 = isu_io_out_valid & exu_io__in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_1 = _T_3 | _GEN_0; // @[Pipeline.scala 26:38]
  reg [63:0] _T_5_cf_instr; // @[Reg.scala 15:16]
  reg [38:0] _T_5_cf_pc; // @[Reg.scala 15:16]
  reg [38:0] _T_5_cf_pnpc; // @[Reg.scala 15:16]
  reg  _T_5_cf_exceptionVec_1; // @[Reg.scala 15:16]
  reg  _T_5_cf_exceptionVec_2; // @[Reg.scala 15:16]
  reg  _T_5_cf_exceptionVec_12; // @[Reg.scala 15:16]
  reg  _T_5_cf_intrVec_0; // @[Reg.scala 15:16]
  reg  _T_5_cf_intrVec_1; // @[Reg.scala 15:16]
  reg  _T_5_cf_intrVec_2; // @[Reg.scala 15:16]
  reg  _T_5_cf_intrVec_3; // @[Reg.scala 15:16]
  reg  _T_5_cf_intrVec_4; // @[Reg.scala 15:16]
  reg  _T_5_cf_intrVec_5; // @[Reg.scala 15:16]
  reg  _T_5_cf_intrVec_6; // @[Reg.scala 15:16]
  reg  _T_5_cf_intrVec_7; // @[Reg.scala 15:16]
  reg  _T_5_cf_intrVec_8; // @[Reg.scala 15:16]
  reg  _T_5_cf_intrVec_9; // @[Reg.scala 15:16]
  reg  _T_5_cf_intrVec_10; // @[Reg.scala 15:16]
  reg  _T_5_cf_intrVec_11; // @[Reg.scala 15:16]
  reg [3:0] _T_5_cf_brIdx; // @[Reg.scala 15:16]
  reg  _T_5_cf_crossPageIPFFix; // @[Reg.scala 15:16]
  reg [2:0] _T_5_ctrl_fuType; // @[Reg.scala 15:16]
  reg [6:0] _T_5_ctrl_fuOpType; // @[Reg.scala 15:16]
  reg  _T_5_ctrl_rfWen; // @[Reg.scala 15:16]
  reg [4:0] _T_5_ctrl_rfDest; // @[Reg.scala 15:16]
  reg [63:0] _T_5_data_src1; // @[Reg.scala 15:16]
  reg [63:0] _T_5_data_src2; // @[Reg.scala 15:16]
  reg [63:0] _T_5_data_imm; // @[Reg.scala 15:16]
  reg  _T_7; // @[Pipeline.scala 24:24]
  wire  _T_8 = exu_io__out_valid; // @[Pipeline.scala 26:22]
  reg [38:0] _T_10_decode_cf_pc; // @[Reg.scala 15:16]
  reg [38:0] _T_10_decode_cf_redirect_target; // @[Reg.scala 15:16]
  reg  _T_10_decode_cf_redirect_valid; // @[Reg.scala 15:16]
  reg [2:0] _T_10_decode_ctrl_fuType; // @[Reg.scala 15:16]
  reg  _T_10_decode_ctrl_rfWen; // @[Reg.scala 15:16]
  reg [4:0] _T_10_decode_ctrl_rfDest; // @[Reg.scala 15:16]
  reg [63:0] _T_10_commits_0; // @[Reg.scala 15:16]
  reg [63:0] _T_10_commits_1; // @[Reg.scala 15:16]
  reg [63:0] _T_10_commits_2; // @[Reg.scala 15:16]
  reg [63:0] _T_10_commits_3; // @[Reg.scala 15:16]
  ISU isu ( // @[Backend.scala 675:20]
    .clock(isu_clock),
    .reset(isu_reset),
    .io_in_0_ready(isu_io_in_0_ready),
    .io_in_0_valid(isu_io_in_0_valid),
    .io_in_0_bits_cf_instr(isu_io_in_0_bits_cf_instr),
    .io_in_0_bits_cf_pc(isu_io_in_0_bits_cf_pc),
    .io_in_0_bits_cf_pnpc(isu_io_in_0_bits_cf_pnpc),
    .io_in_0_bits_cf_exceptionVec_1(isu_io_in_0_bits_cf_exceptionVec_1),
    .io_in_0_bits_cf_exceptionVec_2(isu_io_in_0_bits_cf_exceptionVec_2),
    .io_in_0_bits_cf_exceptionVec_12(isu_io_in_0_bits_cf_exceptionVec_12),
    .io_in_0_bits_cf_intrVec_0(isu_io_in_0_bits_cf_intrVec_0),
    .io_in_0_bits_cf_intrVec_1(isu_io_in_0_bits_cf_intrVec_1),
    .io_in_0_bits_cf_intrVec_2(isu_io_in_0_bits_cf_intrVec_2),
    .io_in_0_bits_cf_intrVec_3(isu_io_in_0_bits_cf_intrVec_3),
    .io_in_0_bits_cf_intrVec_4(isu_io_in_0_bits_cf_intrVec_4),
    .io_in_0_bits_cf_intrVec_5(isu_io_in_0_bits_cf_intrVec_5),
    .io_in_0_bits_cf_intrVec_6(isu_io_in_0_bits_cf_intrVec_6),
    .io_in_0_bits_cf_intrVec_7(isu_io_in_0_bits_cf_intrVec_7),
    .io_in_0_bits_cf_intrVec_8(isu_io_in_0_bits_cf_intrVec_8),
    .io_in_0_bits_cf_intrVec_9(isu_io_in_0_bits_cf_intrVec_9),
    .io_in_0_bits_cf_intrVec_10(isu_io_in_0_bits_cf_intrVec_10),
    .io_in_0_bits_cf_intrVec_11(isu_io_in_0_bits_cf_intrVec_11),
    .io_in_0_bits_cf_brIdx(isu_io_in_0_bits_cf_brIdx),
    .io_in_0_bits_cf_crossPageIPFFix(isu_io_in_0_bits_cf_crossPageIPFFix),
    .io_in_0_bits_ctrl_src1Type(isu_io_in_0_bits_ctrl_src1Type),
    .io_in_0_bits_ctrl_src2Type(isu_io_in_0_bits_ctrl_src2Type),
    .io_in_0_bits_ctrl_fuType(isu_io_in_0_bits_ctrl_fuType),
    .io_in_0_bits_ctrl_fuOpType(isu_io_in_0_bits_ctrl_fuOpType),
    .io_in_0_bits_ctrl_rfSrc1(isu_io_in_0_bits_ctrl_rfSrc1),
    .io_in_0_bits_ctrl_rfSrc2(isu_io_in_0_bits_ctrl_rfSrc2),
    .io_in_0_bits_ctrl_rfWen(isu_io_in_0_bits_ctrl_rfWen),
    .io_in_0_bits_ctrl_rfDest(isu_io_in_0_bits_ctrl_rfDest),
    .io_in_0_bits_data_imm(isu_io_in_0_bits_data_imm),
    .io_out_ready(isu_io_out_ready),
    .io_out_valid(isu_io_out_valid),
    .io_out_bits_cf_instr(isu_io_out_bits_cf_instr),
    .io_out_bits_cf_pc(isu_io_out_bits_cf_pc),
    .io_out_bits_cf_pnpc(isu_io_out_bits_cf_pnpc),
    .io_out_bits_cf_exceptionVec_1(isu_io_out_bits_cf_exceptionVec_1),
    .io_out_bits_cf_exceptionVec_2(isu_io_out_bits_cf_exceptionVec_2),
    .io_out_bits_cf_exceptionVec_12(isu_io_out_bits_cf_exceptionVec_12),
    .io_out_bits_cf_intrVec_0(isu_io_out_bits_cf_intrVec_0),
    .io_out_bits_cf_intrVec_1(isu_io_out_bits_cf_intrVec_1),
    .io_out_bits_cf_intrVec_2(isu_io_out_bits_cf_intrVec_2),
    .io_out_bits_cf_intrVec_3(isu_io_out_bits_cf_intrVec_3),
    .io_out_bits_cf_intrVec_4(isu_io_out_bits_cf_intrVec_4),
    .io_out_bits_cf_intrVec_5(isu_io_out_bits_cf_intrVec_5),
    .io_out_bits_cf_intrVec_6(isu_io_out_bits_cf_intrVec_6),
    .io_out_bits_cf_intrVec_7(isu_io_out_bits_cf_intrVec_7),
    .io_out_bits_cf_intrVec_8(isu_io_out_bits_cf_intrVec_8),
    .io_out_bits_cf_intrVec_9(isu_io_out_bits_cf_intrVec_9),
    .io_out_bits_cf_intrVec_10(isu_io_out_bits_cf_intrVec_10),
    .io_out_bits_cf_intrVec_11(isu_io_out_bits_cf_intrVec_11),
    .io_out_bits_cf_brIdx(isu_io_out_bits_cf_brIdx),
    .io_out_bits_cf_crossPageIPFFix(isu_io_out_bits_cf_crossPageIPFFix),
    .io_out_bits_ctrl_fuType(isu_io_out_bits_ctrl_fuType),
    .io_out_bits_ctrl_fuOpType(isu_io_out_bits_ctrl_fuOpType),
    .io_out_bits_ctrl_rfWen(isu_io_out_bits_ctrl_rfWen),
    .io_out_bits_ctrl_rfDest(isu_io_out_bits_ctrl_rfDest),
    .io_out_bits_data_src1(isu_io_out_bits_data_src1),
    .io_out_bits_data_src2(isu_io_out_bits_data_src2),
    .io_out_bits_data_imm(isu_io_out_bits_data_imm),
    .io_wb_rfWen(isu_io_wb_rfWen),
    .io_wb_rfDest(isu_io_wb_rfDest),
    .io_wb_rfData(isu_io_wb_rfData),
    .io_forward_valid(isu_io_forward_valid),
    .io_forward_wb_rfWen(isu_io_forward_wb_rfWen),
    .io_forward_wb_rfDest(isu_io_forward_wb_rfDest),
    .io_forward_wb_rfData(isu_io_forward_wb_rfData),
    .io_forward_fuType(isu_io_forward_fuType),
    .io_flush(isu_io_flush)
  );
  EXU exu ( // @[Backend.scala 676:20]
    .clock(exu_clock),
    .reset(exu_reset),
    .io__in_ready(exu_io__in_ready),
    .io__in_valid(exu_io__in_valid),
    .io__in_bits_cf_instr(exu_io__in_bits_cf_instr),
    .io__in_bits_cf_pc(exu_io__in_bits_cf_pc),
    .io__in_bits_cf_pnpc(exu_io__in_bits_cf_pnpc),
    .io__in_bits_cf_exceptionVec_1(exu_io__in_bits_cf_exceptionVec_1),
    .io__in_bits_cf_exceptionVec_2(exu_io__in_bits_cf_exceptionVec_2),
    .io__in_bits_cf_exceptionVec_12(exu_io__in_bits_cf_exceptionVec_12),
    .io__in_bits_cf_intrVec_0(exu_io__in_bits_cf_intrVec_0),
    .io__in_bits_cf_intrVec_1(exu_io__in_bits_cf_intrVec_1),
    .io__in_bits_cf_intrVec_2(exu_io__in_bits_cf_intrVec_2),
    .io__in_bits_cf_intrVec_3(exu_io__in_bits_cf_intrVec_3),
    .io__in_bits_cf_intrVec_4(exu_io__in_bits_cf_intrVec_4),
    .io__in_bits_cf_intrVec_5(exu_io__in_bits_cf_intrVec_5),
    .io__in_bits_cf_intrVec_6(exu_io__in_bits_cf_intrVec_6),
    .io__in_bits_cf_intrVec_7(exu_io__in_bits_cf_intrVec_7),
    .io__in_bits_cf_intrVec_8(exu_io__in_bits_cf_intrVec_8),
    .io__in_bits_cf_intrVec_9(exu_io__in_bits_cf_intrVec_9),
    .io__in_bits_cf_intrVec_10(exu_io__in_bits_cf_intrVec_10),
    .io__in_bits_cf_intrVec_11(exu_io__in_bits_cf_intrVec_11),
    .io__in_bits_cf_brIdx(exu_io__in_bits_cf_brIdx),
    .io__in_bits_cf_crossPageIPFFix(exu_io__in_bits_cf_crossPageIPFFix),
    .io__in_bits_ctrl_fuType(exu_io__in_bits_ctrl_fuType),
    .io__in_bits_ctrl_fuOpType(exu_io__in_bits_ctrl_fuOpType),
    .io__in_bits_ctrl_rfWen(exu_io__in_bits_ctrl_rfWen),
    .io__in_bits_ctrl_rfDest(exu_io__in_bits_ctrl_rfDest),
    .io__in_bits_data_src1(exu_io__in_bits_data_src1),
    .io__in_bits_data_src2(exu_io__in_bits_data_src2),
    .io__in_bits_data_imm(exu_io__in_bits_data_imm),
    .io__out_ready(exu_io__out_ready),
    .io__out_valid(exu_io__out_valid),
    .io__out_bits_decode_cf_pc(exu_io__out_bits_decode_cf_pc),
    .io__out_bits_decode_cf_redirect_target(exu_io__out_bits_decode_cf_redirect_target),
    .io__out_bits_decode_cf_redirect_valid(exu_io__out_bits_decode_cf_redirect_valid),
    .io__out_bits_decode_ctrl_fuType(exu_io__out_bits_decode_ctrl_fuType),
    .io__out_bits_decode_ctrl_rfWen(exu_io__out_bits_decode_ctrl_rfWen),
    .io__out_bits_decode_ctrl_rfDest(exu_io__out_bits_decode_ctrl_rfDest),
    .io__out_bits_commits_0(exu_io__out_bits_commits_0),
    .io__out_bits_commits_1(exu_io__out_bits_commits_1),
    .io__out_bits_commits_2(exu_io__out_bits_commits_2),
    .io__out_bits_commits_3(exu_io__out_bits_commits_3),
    .io__flush(exu_io__flush),
    .io__dmem_req_ready(exu_io__dmem_req_ready),
    .io__dmem_req_valid(exu_io__dmem_req_valid),
    .io__dmem_req_bits_addr(exu_io__dmem_req_bits_addr),
    .io__dmem_req_bits_size(exu_io__dmem_req_bits_size),
    .io__dmem_req_bits_cmd(exu_io__dmem_req_bits_cmd),
    .io__dmem_req_bits_wmask(exu_io__dmem_req_bits_wmask),
    .io__dmem_req_bits_wdata(exu_io__dmem_req_bits_wdata),
    .io__dmem_resp_valid(exu_io__dmem_resp_valid),
    .io__dmem_resp_bits_rdata(exu_io__dmem_resp_bits_rdata),
    .io__forward_valid(exu_io__forward_valid),
    .io__forward_wb_rfWen(exu_io__forward_wb_rfWen),
    .io__forward_wb_rfDest(exu_io__forward_wb_rfDest),
    .io__forward_wb_rfData(exu_io__forward_wb_rfData),
    .io__forward_fuType(exu_io__forward_fuType),
    .io__memMMU_imem_priviledgeMode(exu_io__memMMU_imem_priviledgeMode),
    .io__memMMU_dmem_priviledgeMode(exu_io__memMMU_dmem_priviledgeMode),
    .io__memMMU_dmem_status_sum(exu_io__memMMU_dmem_status_sum),
    .io__memMMU_dmem_status_mxr(exu_io__memMMU_dmem_status_mxr),
    .io__memMMU_dmem_loadPF(exu_io__memMMU_dmem_loadPF),
    .io__memMMU_dmem_storePF(exu_io__memMMU_dmem_storePF),
    .io__memMMU_dmem_addr(exu_io__memMMU_dmem_addr),
    ._T_38_0(exu__T_38_0),
    .flushICache(exu_flushICache),
    .perfCnts_2(exu_perfCnts_2),
    .satp(exu_satp),
    ._T_243_valid(exu__T_243_valid),
    ._T_243_pc(exu__T_243_pc),
    ._T_243_isMissPredict(exu__T_243_isMissPredict),
    ._T_243_actualTarget(exu__T_243_actualTarget),
    ._T_243_actualTaken(exu__T_243_actualTaken),
    ._T_243_fuOpType(exu__T_243_fuOpType),
    ._T_243_btbType(exu__T_243_btbType),
    ._T_243_isRVC(exu__T_243_isRVC),
    .io_in_valid(exu_io_in_valid),
    .io_extra_mtip(exu_io_extra_mtip),
    .amoReq(exu_amoReq),
    .io_extra_meip_0(exu_io_extra_meip_0),
    .vmEnable(exu_vmEnable),
    .intrVec(exu_intrVec),
    ._T_37_0(exu__T_37_0),
    .io_extra_msip(exu_io_extra_msip),
    .flushTLB(exu_flushTLB),
    .falseWire(exu_falseWire)
  );
  WBU wbu ( // @[Backend.scala 677:20]
    .io__in_valid(wbu_io__in_valid),
    .io__in_bits_decode_cf_pc(wbu_io__in_bits_decode_cf_pc),
    .io__in_bits_decode_cf_redirect_target(wbu_io__in_bits_decode_cf_redirect_target),
    .io__in_bits_decode_cf_redirect_valid(wbu_io__in_bits_decode_cf_redirect_valid),
    .io__in_bits_decode_ctrl_fuType(wbu_io__in_bits_decode_ctrl_fuType),
    .io__in_bits_decode_ctrl_rfWen(wbu_io__in_bits_decode_ctrl_rfWen),
    .io__in_bits_decode_ctrl_rfDest(wbu_io__in_bits_decode_ctrl_rfDest),
    .io__in_bits_commits_0(wbu_io__in_bits_commits_0),
    .io__in_bits_commits_1(wbu_io__in_bits_commits_1),
    .io__in_bits_commits_2(wbu_io__in_bits_commits_2),
    .io__in_bits_commits_3(wbu_io__in_bits_commits_3),
    .io__wb_rfWen(wbu_io__wb_rfWen),
    .io__wb_rfDest(wbu_io__wb_rfDest),
    .io__wb_rfData(wbu_io__wb_rfData),
    .io__redirect_target(wbu_io__redirect_target),
    .io__redirect_valid(wbu_io__redirect_valid),
    .io_in_bits_decode_cf_pc(wbu_io_in_bits_decode_cf_pc),
    .io_wb_rfDest(wbu_io_wb_rfDest),
    .io_in_valid(wbu_io_in_valid),
    .io_wb_rfWen(wbu_io_wb_rfWen),
    .io_wb_rfData(wbu_io_wb_rfData),
    .io_in_valid_0(wbu_io_in_valid_0),
    .falseWire_0(wbu_falseWire_0)
  );
  assign io_in_0_ready = isu_io_in_0_ready; // @[Backend.scala 682:13]
  assign io_dmem_req_valid = exu_io__dmem_req_valid; // @[Backend.scala 694:11]
  assign io_dmem_req_bits_addr = exu_io__dmem_req_bits_addr; // @[Backend.scala 694:11]
  assign io_dmem_req_bits_size = exu_io__dmem_req_bits_size; // @[Backend.scala 694:11]
  assign io_dmem_req_bits_cmd = exu_io__dmem_req_bits_cmd; // @[Backend.scala 694:11]
  assign io_dmem_req_bits_wmask = exu_io__dmem_req_bits_wmask; // @[Backend.scala 694:11]
  assign io_dmem_req_bits_wdata = exu_io__dmem_req_bits_wdata; // @[Backend.scala 694:11]
  assign io_memMMU_imem_priviledgeMode = exu_io__memMMU_imem_priviledgeMode; // @[Backend.scala 692:18]
  assign io_memMMU_dmem_priviledgeMode = exu_io__memMMU_dmem_priviledgeMode; // @[Backend.scala 693:18]
  assign io_memMMU_dmem_status_sum = exu_io__memMMU_dmem_status_sum; // @[Backend.scala 693:18]
  assign io_memMMU_dmem_status_mxr = exu_io__memMMU_dmem_status_mxr; // @[Backend.scala 693:18]
  assign io_redirect_target = wbu_io__redirect_target; // @[Backend.scala 688:15]
  assign io_redirect_valid = wbu_io__redirect_valid; // @[Backend.scala 688:15]
  assign flushICache = exu_flushICache;
  assign perfCnts_2 = exu_perfCnts_2;
  assign io_in_bits_decode_cf_pc = wbu_io_in_bits_decode_cf_pc;
  assign satp = exu_satp;
  assign _T_243_valid = exu__T_243_valid;
  assign _T_243_pc = exu__T_243_pc;
  assign _T_243_isMissPredict = exu__T_243_isMissPredict;
  assign _T_243_actualTarget = exu__T_243_actualTarget;
  assign _T_243_actualTaken = exu__T_243_actualTaken;
  assign _T_243_fuOpType = exu__T_243_fuOpType;
  assign _T_243_btbType = exu__T_243_btbType;
  assign _T_243_isRVC = exu__T_243_isRVC;
  assign io_wb_rfDest = wbu_io_wb_rfDest;
  assign amoReq = exu_amoReq;
  assign io_wb_rfWen = wbu_io_wb_rfWen;
  assign io_wb_rfData = wbu_io_wb_rfData;
  assign intrVec = exu_intrVec;
  assign flushTLB = exu_flushTLB;
  assign io_in_valid_0 = wbu_io_in_valid_0;
  assign isu_clock = clock;
  assign isu_reset = reset;
  assign isu_io_in_0_valid = io_in_0_valid; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_instr = io_in_0_bits_cf_instr; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_pc = io_in_0_bits_cf_pc; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_pnpc = io_in_0_bits_cf_pnpc; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_exceptionVec_1 = io_in_0_bits_cf_exceptionVec_1; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_exceptionVec_2 = io_in_0_bits_cf_exceptionVec_2; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_exceptionVec_12 = io_in_0_bits_cf_exceptionVec_12; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_intrVec_0 = io_in_0_bits_cf_intrVec_0; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_intrVec_1 = io_in_0_bits_cf_intrVec_1; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_intrVec_2 = io_in_0_bits_cf_intrVec_2; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_intrVec_3 = io_in_0_bits_cf_intrVec_3; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_intrVec_4 = io_in_0_bits_cf_intrVec_4; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_intrVec_5 = io_in_0_bits_cf_intrVec_5; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_intrVec_6 = io_in_0_bits_cf_intrVec_6; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_intrVec_7 = io_in_0_bits_cf_intrVec_7; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_intrVec_8 = io_in_0_bits_cf_intrVec_8; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_intrVec_9 = io_in_0_bits_cf_intrVec_9; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_intrVec_10 = io_in_0_bits_cf_intrVec_10; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_intrVec_11 = io_in_0_bits_cf_intrVec_11; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_brIdx = io_in_0_bits_cf_brIdx; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_cf_crossPageIPFFix = io_in_0_bits_cf_crossPageIPFFix; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_ctrl_src1Type = io_in_0_bits_ctrl_src1Type; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_ctrl_src2Type = io_in_0_bits_ctrl_src2Type; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_ctrl_fuType = io_in_0_bits_ctrl_fuType; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_ctrl_fuOpType = io_in_0_bits_ctrl_fuOpType; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_ctrl_rfSrc1 = io_in_0_bits_ctrl_rfSrc1; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_ctrl_rfSrc2 = io_in_0_bits_ctrl_rfSrc2; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_ctrl_rfWen = io_in_0_bits_ctrl_rfWen; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_ctrl_rfDest = io_in_0_bits_ctrl_rfDest; // @[Backend.scala 682:13]
  assign isu_io_in_0_bits_data_imm = io_in_0_bits_data_imm; // @[Backend.scala 682:13]
  assign isu_io_out_ready = exu_io__in_ready; // @[Pipeline.scala 29:16]
  assign isu_io_wb_rfWen = wbu_io__wb_rfWen; // @[Backend.scala 687:13]
  assign isu_io_wb_rfDest = wbu_io__wb_rfDest; // @[Backend.scala 687:13]
  assign isu_io_wb_rfData = wbu_io__wb_rfData; // @[Backend.scala 687:13]
  assign isu_io_forward_valid = exu_io__forward_valid; // @[Backend.scala 690:18]
  assign isu_io_forward_wb_rfWen = exu_io__forward_wb_rfWen; // @[Backend.scala 690:18]
  assign isu_io_forward_wb_rfDest = exu_io__forward_wb_rfDest; // @[Backend.scala 690:18]
  assign isu_io_forward_wb_rfData = exu_io__forward_wb_rfData; // @[Backend.scala 690:18]
  assign isu_io_forward_fuType = exu_io__forward_fuType; // @[Backend.scala 690:18]
  assign isu_io_flush = io_flush[0]; // @[Backend.scala 684:16]
  assign exu_clock = clock;
  assign exu_reset = reset;
  assign exu_io__in_valid = _T_2; // @[Pipeline.scala 31:17]
  assign exu_io__in_bits_cf_instr = _T_5_cf_instr; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_pc = _T_5_cf_pc; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_pnpc = _T_5_cf_pnpc; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_exceptionVec_1 = _T_5_cf_exceptionVec_1; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_exceptionVec_2 = _T_5_cf_exceptionVec_2; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_exceptionVec_12 = _T_5_cf_exceptionVec_12; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_0 = _T_5_cf_intrVec_0; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_1 = _T_5_cf_intrVec_1; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_2 = _T_5_cf_intrVec_2; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_3 = _T_5_cf_intrVec_3; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_4 = _T_5_cf_intrVec_4; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_5 = _T_5_cf_intrVec_5; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_6 = _T_5_cf_intrVec_6; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_7 = _T_5_cf_intrVec_7; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_8 = _T_5_cf_intrVec_8; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_9 = _T_5_cf_intrVec_9; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_10 = _T_5_cf_intrVec_10; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_intrVec_11 = _T_5_cf_intrVec_11; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_brIdx = _T_5_cf_brIdx; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_cf_crossPageIPFFix = _T_5_cf_crossPageIPFFix; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_fuType = _T_5_ctrl_fuType; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_fuOpType = _T_5_ctrl_fuOpType; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_rfWen = _T_5_ctrl_rfWen; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_ctrl_rfDest = _T_5_ctrl_rfDest; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_data_src1 = _T_5_data_src1; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_data_src2 = _T_5_data_src2; // @[Pipeline.scala 30:16]
  assign exu_io__in_bits_data_imm = _T_5_data_imm; // @[Pipeline.scala 30:16]
  assign exu_io__out_ready = 1'h1; // @[Pipeline.scala 29:16]
  assign exu_io__flush = io_flush[1]; // @[Backend.scala 685:16]
  assign exu_io__dmem_req_ready = io_dmem_req_ready; // @[Backend.scala 694:11]
  assign exu_io__dmem_resp_valid = io_dmem_resp_valid; // @[Backend.scala 694:11]
  assign exu_io__dmem_resp_bits_rdata = io_dmem_resp_bits_rdata; // @[Backend.scala 694:11]
  assign exu_io__memMMU_dmem_loadPF = io_memMMU_dmem_loadPF; // @[Backend.scala 693:18]
  assign exu_io__memMMU_dmem_storePF = io_memMMU_dmem_storePF; // @[Backend.scala 693:18]
  assign exu_io__memMMU_dmem_addr = io_memMMU_dmem_addr; // @[Backend.scala 693:18]
  assign exu__T_38_0 = _T_38;
  assign exu_io_in_valid = wbu_io_in_valid;
  assign exu_io_extra_mtip = io_extra_mtip;
  assign exu_io_extra_meip_0 = io_extra_meip_0;
  assign exu_vmEnable = vmEnable;
  assign exu__T_37_0 = _T_37;
  assign exu_io_extra_msip = io_extra_msip;
  assign exu_falseWire = wbu_falseWire_0;
  assign wbu_io__in_valid = _T_7; // @[Pipeline.scala 31:17]
  assign wbu_io__in_bits_decode_cf_pc = _T_10_decode_cf_pc; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_cf_redirect_target = _T_10_decode_cf_redirect_target; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_cf_redirect_valid = _T_10_decode_cf_redirect_valid; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_fuType = _T_10_decode_ctrl_fuType; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_rfWen = _T_10_decode_ctrl_rfWen; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_decode_ctrl_rfDest = _T_10_decode_ctrl_rfDest; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_0 = _T_10_commits_0; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_1 = _T_10_commits_1; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_2 = _T_10_commits_2; // @[Pipeline.scala 30:16]
  assign wbu_io__in_bits_commits_3 = _T_10_commits_3; // @[Pipeline.scala 30:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_2 = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  _T_5_cf_instr = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  _T_5_cf_pc = _RAND_2[38:0];
  _RAND_3 = {2{`RANDOM}};
  _T_5_cf_pnpc = _RAND_3[38:0];
  _RAND_4 = {1{`RANDOM}};
  _T_5_cf_exceptionVec_1 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_5_cf_exceptionVec_2 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_5_cf_exceptionVec_12 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_5_cf_intrVec_0 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_5_cf_intrVec_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _T_5_cf_intrVec_2 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _T_5_cf_intrVec_3 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_5_cf_intrVec_4 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _T_5_cf_intrVec_5 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _T_5_cf_intrVec_6 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _T_5_cf_intrVec_7 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _T_5_cf_intrVec_8 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  _T_5_cf_intrVec_9 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  _T_5_cf_intrVec_10 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _T_5_cf_intrVec_11 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  _T_5_cf_brIdx = _RAND_19[3:0];
  _RAND_20 = {1{`RANDOM}};
  _T_5_cf_crossPageIPFFix = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _T_5_ctrl_fuType = _RAND_21[2:0];
  _RAND_22 = {1{`RANDOM}};
  _T_5_ctrl_fuOpType = _RAND_22[6:0];
  _RAND_23 = {1{`RANDOM}};
  _T_5_ctrl_rfWen = _RAND_23[0:0];
  _RAND_24 = {1{`RANDOM}};
  _T_5_ctrl_rfDest = _RAND_24[4:0];
  _RAND_25 = {2{`RANDOM}};
  _T_5_data_src1 = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  _T_5_data_src2 = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  _T_5_data_imm = _RAND_27[63:0];
  _RAND_28 = {1{`RANDOM}};
  _T_7 = _RAND_28[0:0];
  _RAND_29 = {2{`RANDOM}};
  _T_10_decode_cf_pc = _RAND_29[38:0];
  _RAND_30 = {2{`RANDOM}};
  _T_10_decode_cf_redirect_target = _RAND_30[38:0];
  _RAND_31 = {1{`RANDOM}};
  _T_10_decode_cf_redirect_valid = _RAND_31[0:0];
  _RAND_32 = {1{`RANDOM}};
  _T_10_decode_ctrl_fuType = _RAND_32[2:0];
  _RAND_33 = {1{`RANDOM}};
  _T_10_decode_ctrl_rfWen = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  _T_10_decode_ctrl_rfDest = _RAND_34[4:0];
  _RAND_35 = {2{`RANDOM}};
  _T_10_commits_0 = _RAND_35[63:0];
  _RAND_36 = {2{`RANDOM}};
  _T_10_commits_1 = _RAND_36[63:0];
  _RAND_37 = {2{`RANDOM}};
  _T_10_commits_2 = _RAND_37[63:0];
  _RAND_38 = {2{`RANDOM}};
  _T_10_commits_3 = _RAND_38[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_2 <= 1'h0;
    end else if (io_flush[0]) begin
      _T_2 <= 1'h0;
    end else begin
      _T_2 <= _GEN_1;
    end
    if (_T_3) begin
      _T_5_cf_instr <= isu_io_out_bits_cf_instr;
    end
    if (_T_3) begin
      _T_5_cf_pc <= isu_io_out_bits_cf_pc;
    end
    if (_T_3) begin
      _T_5_cf_pnpc <= isu_io_out_bits_cf_pnpc;
    end
    if (_T_3) begin
      _T_5_cf_exceptionVec_1 <= isu_io_out_bits_cf_exceptionVec_1;
    end
    if (_T_3) begin
      _T_5_cf_exceptionVec_2 <= isu_io_out_bits_cf_exceptionVec_2;
    end
    if (_T_3) begin
      _T_5_cf_exceptionVec_12 <= isu_io_out_bits_cf_exceptionVec_12;
    end
    if (_T_3) begin
      _T_5_cf_intrVec_0 <= isu_io_out_bits_cf_intrVec_0;
    end
    if (_T_3) begin
      _T_5_cf_intrVec_1 <= isu_io_out_bits_cf_intrVec_1;
    end
    if (_T_3) begin
      _T_5_cf_intrVec_2 <= isu_io_out_bits_cf_intrVec_2;
    end
    if (_T_3) begin
      _T_5_cf_intrVec_3 <= isu_io_out_bits_cf_intrVec_3;
    end
    if (_T_3) begin
      _T_5_cf_intrVec_4 <= isu_io_out_bits_cf_intrVec_4;
    end
    if (_T_3) begin
      _T_5_cf_intrVec_5 <= isu_io_out_bits_cf_intrVec_5;
    end
    if (_T_3) begin
      _T_5_cf_intrVec_6 <= isu_io_out_bits_cf_intrVec_6;
    end
    if (_T_3) begin
      _T_5_cf_intrVec_7 <= isu_io_out_bits_cf_intrVec_7;
    end
    if (_T_3) begin
      _T_5_cf_intrVec_8 <= isu_io_out_bits_cf_intrVec_8;
    end
    if (_T_3) begin
      _T_5_cf_intrVec_9 <= isu_io_out_bits_cf_intrVec_9;
    end
    if (_T_3) begin
      _T_5_cf_intrVec_10 <= isu_io_out_bits_cf_intrVec_10;
    end
    if (_T_3) begin
      _T_5_cf_intrVec_11 <= isu_io_out_bits_cf_intrVec_11;
    end
    if (_T_3) begin
      _T_5_cf_brIdx <= isu_io_out_bits_cf_brIdx;
    end
    if (_T_3) begin
      _T_5_cf_crossPageIPFFix <= isu_io_out_bits_cf_crossPageIPFFix;
    end
    if (_T_3) begin
      _T_5_ctrl_fuType <= isu_io_out_bits_ctrl_fuType;
    end
    if (_T_3) begin
      _T_5_ctrl_fuOpType <= isu_io_out_bits_ctrl_fuOpType;
    end
    if (_T_3) begin
      _T_5_ctrl_rfWen <= isu_io_out_bits_ctrl_rfWen;
    end
    if (_T_3) begin
      _T_5_ctrl_rfDest <= isu_io_out_bits_ctrl_rfDest;
    end
    if (_T_3) begin
      _T_5_data_src1 <= isu_io_out_bits_data_src1;
    end
    if (_T_3) begin
      _T_5_data_src2 <= isu_io_out_bits_data_src2;
    end
    if (_T_3) begin
      _T_5_data_imm <= isu_io_out_bits_data_imm;
    end
    if (reset) begin
      _T_7 <= 1'h0;
    end else if (io_flush[1]) begin
      _T_7 <= 1'h0;
    end else begin
      _T_7 <= _T_8;
    end
    if (_T_8) begin
      _T_10_decode_cf_pc <= exu_io__out_bits_decode_cf_pc;
    end
    if (_T_8) begin
      _T_10_decode_cf_redirect_target <= exu_io__out_bits_decode_cf_redirect_target;
    end
    if (_T_8) begin
      _T_10_decode_cf_redirect_valid <= exu_io__out_bits_decode_cf_redirect_valid;
    end
    if (_T_8) begin
      _T_10_decode_ctrl_fuType <= exu_io__out_bits_decode_ctrl_fuType;
    end
    if (_T_8) begin
      _T_10_decode_ctrl_rfWen <= exu_io__out_bits_decode_ctrl_rfWen;
    end
    if (_T_8) begin
      _T_10_decode_ctrl_rfDest <= exu_io__out_bits_decode_ctrl_rfDest;
    end
    if (_T_8) begin
      _T_10_commits_0 <= exu_io__out_bits_commits_0;
    end
    if (_T_8) begin
      _T_10_commits_1 <= exu_io__out_bits_commits_1;
    end
    if (_T_8) begin
      _T_10_commits_2 <= exu_io__out_bits_commits_2;
    end
    if (_T_8) begin
      _T_10_commits_3 <= exu_io__out_bits_commits_3;
    end
  end
endmodule
module LockingArbiter(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [3:0]  io_in_0_bits_cmd,
  input  [7:0]  io_in_0_bits_wmask,
  input  [63:0] io_in_0_bits_wdata,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [2:0]  io_in_1_bits_size,
  input  [3:0]  io_in_1_bits_cmd,
  input  [7:0]  io_in_1_bits_wmask,
  input  [63:0] io_in_1_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [2:0]  io_out_bits_size,
  output [3:0]  io_out_bits_cmd,
  output [7:0]  io_out_bits_wmask,
  output [63:0] io_out_bits_wdata,
  output        io_chosen
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] value; // @[Counter.scala 29:33]
  reg  _T; // @[Arbiter.scala 46:22]
  wire  _T_1 = value != 3'h0; // @[Arbiter.scala 47:34]
  wire  _T_4 = io_out_bits_cmd[0] & io_out_bits_cmd[1]; // @[Crossbar.scala 100:62]
  wire  _T_5 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_6 = _T_5 & _T_4; // @[Arbiter.scala 50:25]
  wire [2:0] _T_9 = value + 3'h1; // @[Counter.scala 39:22]
  wire  choice = io_in_0_valid ? 1'h0 : 1'h1; // @[Arbiter.scala 88:27]
  wire  _T_10 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  _T_11 = ~_T; // @[Arbiter.scala 57:39]
  wire  _T_12 = _T_1 ? _T_11 : 1'h1; // @[Arbiter.scala 57:22]
  wire  _T_15 = _T_1 ? _T : _T_10; // @[Arbiter.scala 57:22]
  assign io_in_0_ready = _T_12 & io_out_ready; // @[Arbiter.scala 57:16]
  assign io_in_1_ready = _T_15 & io_out_ready; // @[Arbiter.scala 57:16]
  assign io_out_valid = io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:16]
  assign io_out_bits_addr = io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[Arbiter.scala 42:15]
  assign io_out_bits_size = io_chosen ? io_in_1_bits_size : 3'h3; // @[Arbiter.scala 42:15]
  assign io_out_bits_cmd = io_chosen ? io_in_1_bits_cmd : io_in_0_bits_cmd; // @[Arbiter.scala 42:15]
  assign io_out_bits_wmask = io_chosen ? io_in_1_bits_wmask : io_in_0_bits_wmask; // @[Arbiter.scala 42:15]
  assign io_out_bits_wdata = io_chosen ? io_in_1_bits_wdata : io_in_0_bits_wdata; // @[Arbiter.scala 42:15]
  assign io_chosen = _T_1 ? _T : choice; // @[Arbiter.scala 40:13 Arbiter.scala 55:31]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  _T = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 3'h0;
    end else if (_T_6) begin
      value <= _T_9;
    end
    if (_T_6) begin
      _T <= io_chosen;
    end
  end
endmodule
module SimpleBusCrossbarNto1(
  input         clock,
  input         reset,
  output        io_in_0_req_ready,
  input         io_in_0_req_valid,
  input  [31:0] io_in_0_req_bits_addr,
  input  [3:0]  io_in_0_req_bits_cmd,
  input  [7:0]  io_in_0_req_bits_wmask,
  input  [63:0] io_in_0_req_bits_wdata,
  output        io_in_0_resp_valid,
  output [3:0]  io_in_0_resp_bits_cmd,
  output [63:0] io_in_0_resp_bits_rdata,
  output        io_in_1_req_ready,
  input         io_in_1_req_valid,
  input  [31:0] io_in_1_req_bits_addr,
  input  [2:0]  io_in_1_req_bits_size,
  input  [3:0]  io_in_1_req_bits_cmd,
  input  [7:0]  io_in_1_req_bits_wmask,
  input  [63:0] io_in_1_req_bits_wdata,
  output        io_in_1_resp_valid,
  output [3:0]  io_in_1_resp_bits_cmd,
  output [63:0] io_in_1_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [2:0]  io_out_req_bits_size,
  output [3:0]  io_out_req_bits_cmd,
  output [7:0]  io_out_req_bits_wmask,
  output [63:0] io_out_req_bits_wdata,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [3:0]  io_out_resp_bits_cmd,
  input  [63:0] io_out_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  inputArb_clock; // @[Crossbar.scala 101:24]
  wire  inputArb_reset; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_0_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_0_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_in_0_bits_addr; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_in_0_bits_cmd; // @[Crossbar.scala 101:24]
  wire [7:0] inputArb_io_in_0_bits_wmask; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_in_0_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_1_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_1_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_in_1_bits_addr; // @[Crossbar.scala 101:24]
  wire [2:0] inputArb_io_in_1_bits_size; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_in_1_bits_cmd; // @[Crossbar.scala 101:24]
  wire [7:0] inputArb_io_in_1_bits_wmask; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_in_1_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_out_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_out_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_out_bits_addr; // @[Crossbar.scala 101:24]
  wire [2:0] inputArb_io_out_bits_size; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_out_bits_cmd; // @[Crossbar.scala 101:24]
  wire [7:0] inputArb_io_out_bits_wmask; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_out_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_chosen; // @[Crossbar.scala 101:24]
  reg [1:0] state; // @[Crossbar.scala 98:22]
  wire  _T_1 = ~inputArb_io_out_bits_cmd[0]; // @[SimpleBus.scala 73:18]
  wire  _T_3 = ~inputArb_io_out_bits_cmd[3]; // @[SimpleBus.scala 73:29]
  wire  _T_4 = _T_1 & _T_3; // @[SimpleBus.scala 73:26]
  wire  _T_5 = ~_T_4; // @[Crossbar.scala 104:29]
  wire  _T_6 = inputArb_io_out_valid & _T_5; // @[Crossbar.scala 104:26]
  wire  _T_9 = _T_6 & _T_1; // @[Crossbar.scala 104:52]
  wire  _T_10 = ~_T_9; // @[Crossbar.scala 104:10]
  wire  _T_12 = _T_10 | reset; // @[Crossbar.scala 104:9]
  wire  _T_13 = ~_T_12; // @[Crossbar.scala 104:9]
  reg  inflightSrc; // @[Crossbar.scala 105:24]
  wire  _T_14 = state == 2'h0; // @[Crossbar.scala 109:47]
  wire  _GEN_34 = ~inflightSrc; // @[Crossbar.scala 115:13]
  wire  _T_18 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_19 = inputArb_io_out_ready & inputArb_io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_25 = inputArb_io_out_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_26 = inputArb_io_out_bits_cmd == 4'h1; // @[SimpleBus.scala 77:29]
  wire  _T_27 = _T_25 | _T_26; // @[Crossbar.scala 124:47]
  wire  _T_28 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_29 = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_30 = io_out_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire  _T_31 = _T_29 & _T_30; // @[Crossbar.scala 127:48]
  wire  _T_32 = 2'h2 == state; // @[Conditional.scala 37:30]
  LockingArbiter inputArb ( // @[Crossbar.scala 101:24]
    .clock(inputArb_clock),
    .reset(inputArb_reset),
    .io_in_0_ready(inputArb_io_in_0_ready),
    .io_in_0_valid(inputArb_io_in_0_valid),
    .io_in_0_bits_addr(inputArb_io_in_0_bits_addr),
    .io_in_0_bits_cmd(inputArb_io_in_0_bits_cmd),
    .io_in_0_bits_wmask(inputArb_io_in_0_bits_wmask),
    .io_in_0_bits_wdata(inputArb_io_in_0_bits_wdata),
    .io_in_1_ready(inputArb_io_in_1_ready),
    .io_in_1_valid(inputArb_io_in_1_valid),
    .io_in_1_bits_addr(inputArb_io_in_1_bits_addr),
    .io_in_1_bits_size(inputArb_io_in_1_bits_size),
    .io_in_1_bits_cmd(inputArb_io_in_1_bits_cmd),
    .io_in_1_bits_wmask(inputArb_io_in_1_bits_wmask),
    .io_in_1_bits_wdata(inputArb_io_in_1_bits_wdata),
    .io_out_ready(inputArb_io_out_ready),
    .io_out_valid(inputArb_io_out_valid),
    .io_out_bits_addr(inputArb_io_out_bits_addr),
    .io_out_bits_size(inputArb_io_out_bits_size),
    .io_out_bits_cmd(inputArb_io_out_bits_cmd),
    .io_out_bits_wmask(inputArb_io_out_bits_wmask),
    .io_out_bits_wdata(inputArb_io_out_bits_wdata),
    .io_chosen(inputArb_io_chosen)
  );
  assign io_in_0_req_ready = inputArb_io_in_0_ready; // @[Crossbar.scala 102:68]
  assign io_in_0_resp_valid = _GEN_34 & io_out_resp_valid; // @[Crossbar.scala 113:26 Crossbar.scala 115:13]
  assign io_in_0_resp_bits_cmd = io_out_resp_bits_cmd; // @[Crossbar.scala 112:25]
  assign io_in_0_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 112:25]
  assign io_in_1_req_ready = inputArb_io_in_1_ready; // @[Crossbar.scala 102:68]
  assign io_in_1_resp_valid = inflightSrc & io_out_resp_valid; // @[Crossbar.scala 113:26 Crossbar.scala 115:13]
  assign io_in_1_resp_bits_cmd = io_out_resp_bits_cmd; // @[Crossbar.scala 112:25]
  assign io_in_1_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 112:25]
  assign io_out_req_valid = inputArb_io_out_valid & _T_14; // @[Crossbar.scala 109:20]
  assign io_out_req_bits_addr = inputArb_io_out_bits_addr; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_size = inputArb_io_out_bits_size; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_cmd = inputArb_io_out_bits_cmd; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_wmask = inputArb_io_out_bits_wmask; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_wdata = inputArb_io_out_bits_wdata; // @[Crossbar.scala 107:19]
  assign io_out_resp_ready = 1'h1; // @[Crossbar.scala 116:13]
  assign inputArb_clock = clock;
  assign inputArb_reset = reset;
  assign inputArb_io_in_0_valid = io_in_0_req_valid; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_addr = io_in_0_req_bits_addr; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_cmd = io_in_0_req_bits_cmd; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_wmask = io_in_0_req_bits_wmask; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_wdata = io_in_0_req_bits_wdata; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_valid = io_in_1_req_valid; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_addr = io_in_1_req_bits_addr; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_size = io_in_1_req_bits_size; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_cmd = io_in_1_req_bits_cmd; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_wmask = io_in_1_req_bits_wmask; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_wdata = io_in_1_req_bits_wdata; // @[Crossbar.scala 102:68]
  assign inputArb_io_out_ready = io_out_req_ready & _T_14; // @[Crossbar.scala 110:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  inflightSrc = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else if (_T_18) begin
      if (_T_19) begin
        if (_T_4) begin
          state <= 2'h1;
        end else if (_T_27) begin
          state <= 2'h2;
        end
      end
    end else if (_T_28) begin
      if (_T_31) begin
        state <= 2'h0;
      end
    end else if (_T_32) begin
      if (_T_29) begin
        state <= 2'h0;
      end
    end
    if (_T_18) begin
      if (_T_19) begin
        inflightSrc <= inputArb_io_chosen;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Crossbar.scala:104 assert(!(thisReq.valid && !thisReq.bits.isRead() && !thisReq.bits.isWrite()))\n"); // @[Crossbar.scala 104:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_13) begin
          $fatal; // @[Crossbar.scala 104:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module LockingArbiter_1(
  input         clock,
  input         reset,
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [2:0]  io_in_0_bits_size,
  input  [3:0]  io_in_0_bits_cmd,
  input  [7:0]  io_in_0_bits_wmask,
  input  [63:0] io_in_0_bits_wdata,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [3:0]  io_in_1_bits_cmd,
  input  [63:0] io_in_1_bits_wdata,
  output        io_in_2_ready,
  input         io_in_2_valid,
  input  [31:0] io_in_2_bits_addr,
  input  [3:0]  io_in_2_bits_cmd,
  input  [63:0] io_in_2_bits_wdata,
  output        io_in_3_ready,
  input         io_in_3_valid,
  input  [31:0] io_in_3_bits_addr,
  input  [2:0]  io_in_3_bits_size,
  input  [3:0]  io_in_3_bits_cmd,
  input  [7:0]  io_in_3_bits_wmask,
  input  [63:0] io_in_3_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [2:0]  io_out_bits_size,
  output [3:0]  io_out_bits_cmd,
  output [7:0]  io_out_bits_wmask,
  output [63:0] io_out_bits_wdata,
  output [1:0]  io_chosen
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  _GEN_8 = 2'h1 == io_chosen ? io_in_1_valid : io_in_0_valid; // @[Arbiter.scala 41:16]
  wire [31:0] _GEN_9 = 2'h1 == io_chosen ? io_in_1_bits_addr : io_in_0_bits_addr; // @[Arbiter.scala 41:16]
  wire [2:0] _GEN_10 = 2'h1 == io_chosen ? 3'h3 : io_in_0_bits_size; // @[Arbiter.scala 41:16]
  wire [3:0] _GEN_11 = 2'h1 == io_chosen ? io_in_1_bits_cmd : io_in_0_bits_cmd; // @[Arbiter.scala 41:16]
  wire [7:0] _GEN_12 = 2'h1 == io_chosen ? 8'hff : io_in_0_bits_wmask; // @[Arbiter.scala 41:16]
  wire [63:0] _GEN_13 = 2'h1 == io_chosen ? io_in_1_bits_wdata : io_in_0_bits_wdata; // @[Arbiter.scala 41:16]
  wire  _GEN_15 = 2'h2 == io_chosen ? io_in_2_valid : _GEN_8; // @[Arbiter.scala 41:16]
  wire [31:0] _GEN_16 = 2'h2 == io_chosen ? io_in_2_bits_addr : _GEN_9; // @[Arbiter.scala 41:16]
  wire [2:0] _GEN_17 = 2'h2 == io_chosen ? 3'h3 : _GEN_10; // @[Arbiter.scala 41:16]
  wire [3:0] _GEN_18 = 2'h2 == io_chosen ? io_in_2_bits_cmd : _GEN_11; // @[Arbiter.scala 41:16]
  wire [7:0] _GEN_19 = 2'h2 == io_chosen ? 8'hff : _GEN_12; // @[Arbiter.scala 41:16]
  wire [63:0] _GEN_20 = 2'h2 == io_chosen ? io_in_2_bits_wdata : _GEN_13; // @[Arbiter.scala 41:16]
  reg [2:0] value; // @[Counter.scala 29:33]
  reg [1:0] _T; // @[Arbiter.scala 46:22]
  wire  _T_1 = value != 3'h0; // @[Arbiter.scala 47:34]
  wire  _T_4 = io_out_bits_cmd[0] & io_out_bits_cmd[1]; // @[Crossbar.scala 100:62]
  wire  _T_5 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_6 = _T_5 & _T_4; // @[Arbiter.scala 50:25]
  wire [2:0] _T_9 = value + 3'h1; // @[Counter.scala 39:22]
  wire [1:0] _GEN_31 = io_in_2_valid ? 2'h2 : 2'h3; // @[Arbiter.scala 88:27]
  wire [1:0] _GEN_32 = io_in_1_valid ? 2'h1 : _GEN_31; // @[Arbiter.scala 88:27]
  wire [1:0] choice = io_in_0_valid ? 2'h0 : _GEN_32; // @[Arbiter.scala 88:27]
  wire  _T_10 = io_in_0_valid | io_in_1_valid; // @[Arbiter.scala 31:68]
  wire  _T_11 = _T_10 | io_in_2_valid; // @[Arbiter.scala 31:68]
  wire  _T_12 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  _T_13 = ~_T_10; // @[Arbiter.scala 31:78]
  wire  _T_14 = ~_T_11; // @[Arbiter.scala 31:78]
  wire  _T_15 = _T == 2'h0; // @[Arbiter.scala 57:39]
  wire  _T_16 = _T_1 ? _T_15 : 1'h1; // @[Arbiter.scala 57:22]
  wire  _T_18 = _T == 2'h1; // @[Arbiter.scala 57:39]
  wire  _T_19 = _T_1 ? _T_18 : _T_12; // @[Arbiter.scala 57:22]
  wire  _T_21 = _T == 2'h2; // @[Arbiter.scala 57:39]
  wire  _T_22 = _T_1 ? _T_21 : _T_13; // @[Arbiter.scala 57:22]
  wire  _T_24 = _T == 2'h3; // @[Arbiter.scala 57:39]
  wire  _T_25 = _T_1 ? _T_24 : _T_14; // @[Arbiter.scala 57:22]
  assign io_in_0_ready = _T_16 & io_out_ready; // @[Arbiter.scala 57:16]
  assign io_in_1_ready = _T_19 & io_out_ready; // @[Arbiter.scala 57:16]
  assign io_in_2_ready = _T_22 & io_out_ready; // @[Arbiter.scala 57:16]
  assign io_in_3_ready = _T_25 & io_out_ready; // @[Arbiter.scala 57:16]
  assign io_out_valid = 2'h3 == io_chosen ? io_in_3_valid : _GEN_15; // @[Arbiter.scala 41:16]
  assign io_out_bits_addr = 2'h3 == io_chosen ? io_in_3_bits_addr : _GEN_16; // @[Arbiter.scala 42:15]
  assign io_out_bits_size = 2'h3 == io_chosen ? io_in_3_bits_size : _GEN_17; // @[Arbiter.scala 42:15]
  assign io_out_bits_cmd = 2'h3 == io_chosen ? io_in_3_bits_cmd : _GEN_18; // @[Arbiter.scala 42:15]
  assign io_out_bits_wmask = 2'h3 == io_chosen ? io_in_3_bits_wmask : _GEN_19; // @[Arbiter.scala 42:15]
  assign io_out_bits_wdata = 2'h3 == io_chosen ? io_in_3_bits_wdata : _GEN_20; // @[Arbiter.scala 42:15]
  assign io_chosen = _T_1 ? _T : choice; // @[Arbiter.scala 40:13 Arbiter.scala 55:31]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  _T = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 3'h0;
    end else if (_T_6) begin
      value <= _T_9;
    end
    if (_T_6) begin
      _T <= io_chosen;
    end
  end
endmodule
module SimpleBusCrossbarNto1_1(
  input         clock,
  input         reset,
  output        io_in_0_req_ready,
  input         io_in_0_req_valid,
  input  [31:0] io_in_0_req_bits_addr,
  input  [2:0]  io_in_0_req_bits_size,
  input  [3:0]  io_in_0_req_bits_cmd,
  input  [7:0]  io_in_0_req_bits_wmask,
  input  [63:0] io_in_0_req_bits_wdata,
  output        io_in_0_resp_valid,
  output [63:0] io_in_0_resp_bits_rdata,
  output        io_in_1_req_ready,
  input         io_in_1_req_valid,
  input  [31:0] io_in_1_req_bits_addr,
  input  [3:0]  io_in_1_req_bits_cmd,
  input  [63:0] io_in_1_req_bits_wdata,
  output        io_in_1_resp_valid,
  output [63:0] io_in_1_resp_bits_rdata,
  output        io_in_2_req_ready,
  input         io_in_2_req_valid,
  input  [31:0] io_in_2_req_bits_addr,
  input  [3:0]  io_in_2_req_bits_cmd,
  input  [63:0] io_in_2_req_bits_wdata,
  output        io_in_2_resp_valid,
  output [63:0] io_in_2_resp_bits_rdata,
  output        io_in_3_req_ready,
  input         io_in_3_req_valid,
  input  [31:0] io_in_3_req_bits_addr,
  input  [2:0]  io_in_3_req_bits_size,
  input  [3:0]  io_in_3_req_bits_cmd,
  input  [7:0]  io_in_3_req_bits_wmask,
  input  [63:0] io_in_3_req_bits_wdata,
  input         io_in_3_resp_ready,
  output        io_in_3_resp_valid,
  output [3:0]  io_in_3_resp_bits_cmd,
  output [63:0] io_in_3_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [2:0]  io_out_req_bits_size,
  output [3:0]  io_out_req_bits_cmd,
  output [7:0]  io_out_req_bits_wmask,
  output [63:0] io_out_req_bits_wdata,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [3:0]  io_out_resp_bits_cmd,
  input  [63:0] io_out_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  inputArb_clock; // @[Crossbar.scala 101:24]
  wire  inputArb_reset; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_0_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_0_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_in_0_bits_addr; // @[Crossbar.scala 101:24]
  wire [2:0] inputArb_io_in_0_bits_size; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_in_0_bits_cmd; // @[Crossbar.scala 101:24]
  wire [7:0] inputArb_io_in_0_bits_wmask; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_in_0_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_1_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_1_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_in_1_bits_addr; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_in_1_bits_cmd; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_in_1_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_2_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_2_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_in_2_bits_addr; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_in_2_bits_cmd; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_in_2_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_3_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_in_3_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_in_3_bits_addr; // @[Crossbar.scala 101:24]
  wire [2:0] inputArb_io_in_3_bits_size; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_in_3_bits_cmd; // @[Crossbar.scala 101:24]
  wire [7:0] inputArb_io_in_3_bits_wmask; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_in_3_bits_wdata; // @[Crossbar.scala 101:24]
  wire  inputArb_io_out_ready; // @[Crossbar.scala 101:24]
  wire  inputArb_io_out_valid; // @[Crossbar.scala 101:24]
  wire [31:0] inputArb_io_out_bits_addr; // @[Crossbar.scala 101:24]
  wire [2:0] inputArb_io_out_bits_size; // @[Crossbar.scala 101:24]
  wire [3:0] inputArb_io_out_bits_cmd; // @[Crossbar.scala 101:24]
  wire [7:0] inputArb_io_out_bits_wmask; // @[Crossbar.scala 101:24]
  wire [63:0] inputArb_io_out_bits_wdata; // @[Crossbar.scala 101:24]
  wire [1:0] inputArb_io_chosen; // @[Crossbar.scala 101:24]
  reg [1:0] state; // @[Crossbar.scala 98:22]
  wire  _T_1 = ~inputArb_io_out_bits_cmd[0]; // @[SimpleBus.scala 73:18]
  wire  _T_3 = ~inputArb_io_out_bits_cmd[3]; // @[SimpleBus.scala 73:29]
  wire  _T_4 = _T_1 & _T_3; // @[SimpleBus.scala 73:26]
  wire  _T_5 = ~_T_4; // @[Crossbar.scala 104:29]
  wire  _T_6 = inputArb_io_out_valid & _T_5; // @[Crossbar.scala 104:26]
  wire  _T_9 = _T_6 & _T_1; // @[Crossbar.scala 104:52]
  wire  _T_10 = ~_T_9; // @[Crossbar.scala 104:10]
  wire  _T_12 = _T_10 | reset; // @[Crossbar.scala 104:9]
  wire  _T_13 = ~_T_12; // @[Crossbar.scala 104:9]
  reg [1:0] inflightSrc; // @[Crossbar.scala 105:24]
  wire  _T_14 = state == 2'h0; // @[Crossbar.scala 109:47]
  wire  _GEN_58 = 2'h0 == inflightSrc; // @[Crossbar.scala 115:13]
  wire  _GEN_59 = 2'h1 == inflightSrc; // @[Crossbar.scala 115:13]
  wire  _GEN_60 = 2'h2 == inflightSrc; // @[Crossbar.scala 115:13]
  wire  _GEN_61 = 2'h3 == inflightSrc; // @[Crossbar.scala 115:13]
  wire  _T_18 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_19 = inputArb_io_out_ready & inputArb_io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_25 = inputArb_io_out_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_26 = inputArb_io_out_bits_cmd == 4'h1; // @[SimpleBus.scala 77:29]
  wire  _T_27 = _T_25 | _T_26; // @[Crossbar.scala 124:47]
  wire  _T_28 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_29 = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_30 = io_out_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire  _T_31 = _T_29 & _T_30; // @[Crossbar.scala 127:48]
  wire  _T_32 = 2'h2 == state; // @[Conditional.scala 37:30]
  LockingArbiter_1 inputArb ( // @[Crossbar.scala 101:24]
    .clock(inputArb_clock),
    .reset(inputArb_reset),
    .io_in_0_ready(inputArb_io_in_0_ready),
    .io_in_0_valid(inputArb_io_in_0_valid),
    .io_in_0_bits_addr(inputArb_io_in_0_bits_addr),
    .io_in_0_bits_size(inputArb_io_in_0_bits_size),
    .io_in_0_bits_cmd(inputArb_io_in_0_bits_cmd),
    .io_in_0_bits_wmask(inputArb_io_in_0_bits_wmask),
    .io_in_0_bits_wdata(inputArb_io_in_0_bits_wdata),
    .io_in_1_ready(inputArb_io_in_1_ready),
    .io_in_1_valid(inputArb_io_in_1_valid),
    .io_in_1_bits_addr(inputArb_io_in_1_bits_addr),
    .io_in_1_bits_cmd(inputArb_io_in_1_bits_cmd),
    .io_in_1_bits_wdata(inputArb_io_in_1_bits_wdata),
    .io_in_2_ready(inputArb_io_in_2_ready),
    .io_in_2_valid(inputArb_io_in_2_valid),
    .io_in_2_bits_addr(inputArb_io_in_2_bits_addr),
    .io_in_2_bits_cmd(inputArb_io_in_2_bits_cmd),
    .io_in_2_bits_wdata(inputArb_io_in_2_bits_wdata),
    .io_in_3_ready(inputArb_io_in_3_ready),
    .io_in_3_valid(inputArb_io_in_3_valid),
    .io_in_3_bits_addr(inputArb_io_in_3_bits_addr),
    .io_in_3_bits_size(inputArb_io_in_3_bits_size),
    .io_in_3_bits_cmd(inputArb_io_in_3_bits_cmd),
    .io_in_3_bits_wmask(inputArb_io_in_3_bits_wmask),
    .io_in_3_bits_wdata(inputArb_io_in_3_bits_wdata),
    .io_out_ready(inputArb_io_out_ready),
    .io_out_valid(inputArb_io_out_valid),
    .io_out_bits_addr(inputArb_io_out_bits_addr),
    .io_out_bits_size(inputArb_io_out_bits_size),
    .io_out_bits_cmd(inputArb_io_out_bits_cmd),
    .io_out_bits_wmask(inputArb_io_out_bits_wmask),
    .io_out_bits_wdata(inputArb_io_out_bits_wdata),
    .io_chosen(inputArb_io_chosen)
  );
  assign io_in_0_req_ready = inputArb_io_in_0_ready; // @[Crossbar.scala 102:68]
  assign io_in_0_resp_valid = _GEN_58 & io_out_resp_valid; // @[Crossbar.scala 113:26 Crossbar.scala 115:13]
  assign io_in_0_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 112:25]
  assign io_in_1_req_ready = inputArb_io_in_1_ready; // @[Crossbar.scala 102:68]
  assign io_in_1_resp_valid = _GEN_59 & io_out_resp_valid; // @[Crossbar.scala 113:26 Crossbar.scala 115:13]
  assign io_in_1_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 112:25]
  assign io_in_2_req_ready = inputArb_io_in_2_ready; // @[Crossbar.scala 102:68]
  assign io_in_2_resp_valid = _GEN_60 & io_out_resp_valid; // @[Crossbar.scala 113:26 Crossbar.scala 115:13]
  assign io_in_2_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 112:25]
  assign io_in_3_req_ready = inputArb_io_in_3_ready; // @[Crossbar.scala 102:68]
  assign io_in_3_resp_valid = _GEN_61 & io_out_resp_valid; // @[Crossbar.scala 113:26 Crossbar.scala 115:13]
  assign io_in_3_resp_bits_cmd = io_out_resp_bits_cmd; // @[Crossbar.scala 112:25]
  assign io_in_3_resp_bits_rdata = io_out_resp_bits_rdata; // @[Crossbar.scala 112:25]
  assign io_out_req_valid = inputArb_io_out_valid & _T_14; // @[Crossbar.scala 109:20]
  assign io_out_req_bits_addr = inputArb_io_out_bits_addr; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_size = inputArb_io_out_bits_size; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_cmd = inputArb_io_out_bits_cmd; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_wmask = inputArb_io_out_bits_wmask; // @[Crossbar.scala 107:19]
  assign io_out_req_bits_wdata = inputArb_io_out_bits_wdata; // @[Crossbar.scala 107:19]
  assign io_out_resp_ready = 2'h3 == inflightSrc ? io_in_3_resp_ready : 1'h1; // @[Crossbar.scala 116:13]
  assign inputArb_clock = clock;
  assign inputArb_reset = reset;
  assign inputArb_io_in_0_valid = io_in_0_req_valid; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_addr = io_in_0_req_bits_addr; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_size = io_in_0_req_bits_size; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_cmd = io_in_0_req_bits_cmd; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_wmask = io_in_0_req_bits_wmask; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_0_bits_wdata = io_in_0_req_bits_wdata; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_valid = io_in_1_req_valid; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_addr = io_in_1_req_bits_addr; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_cmd = io_in_1_req_bits_cmd; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_1_bits_wdata = io_in_1_req_bits_wdata; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_2_valid = io_in_2_req_valid; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_2_bits_addr = io_in_2_req_bits_addr; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_2_bits_cmd = io_in_2_req_bits_cmd; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_2_bits_wdata = io_in_2_req_bits_wdata; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_3_valid = io_in_3_req_valid; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_3_bits_addr = io_in_3_req_bits_addr; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_3_bits_size = io_in_3_req_bits_size; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_3_bits_cmd = io_in_3_req_bits_cmd; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_3_bits_wmask = io_in_3_req_bits_wmask; // @[Crossbar.scala 102:68]
  assign inputArb_io_in_3_bits_wdata = io_in_3_req_bits_wdata; // @[Crossbar.scala 102:68]
  assign inputArb_io_out_ready = io_out_req_ready & _T_14; // @[Crossbar.scala 110:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  inflightSrc = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else if (_T_18) begin
      if (_T_19) begin
        if (_T_4) begin
          state <= 2'h1;
        end else if (_T_27) begin
          state <= 2'h2;
        end
      end
    end else if (_T_28) begin
      if (_T_31) begin
        state <= 2'h0;
      end
    end else if (_T_32) begin
      if (_T_29) begin
        state <= 2'h0;
      end
    end
    if (_T_18) begin
      if (_T_19) begin
        inflightSrc <= inputArb_io_chosen;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Crossbar.scala:104 assert(!(thisReq.valid && !thisReq.bits.isRead() && !thisReq.bits.isWrite()))\n"); // @[Crossbar.scala 104:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_13) begin
          $fatal; // @[Crossbar.scala 104:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module EmbeddedTLBExec(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [38:0]  io_in_bits_addr,
  input  [86:0]  io_in_bits_user,
  input          io_out_ready,
  output         io_out_valid,
  output [31:0]  io_out_bits_addr,
  output [86:0]  io_out_bits_user,
  input  [120:0] io_md_0,
  input  [120:0] io_md_1,
  input  [120:0] io_md_2,
  input  [120:0] io_md_3,
  output         io_mdWrite_wen,
  output [3:0]   io_mdWrite_waymask,
  output [120:0] io_mdWrite_wdata,
  input          io_mdReady,
  input          io_mem_req_ready,
  output         io_mem_req_valid,
  output [31:0]  io_mem_req_bits_addr,
  output [3:0]   io_mem_req_bits_cmd,
  output [63:0]  io_mem_req_bits_wdata,
  output         io_mem_resp_ready,
  input          io_mem_resp_valid,
  input  [63:0]  io_mem_resp_bits_rdata,
  input          io_flush,
  input  [63:0]  io_satp,
  input  [1:0]   io_pf_priviledgeMode,
  output         io_pf_loadPF,
  output         io_pf_storePF,
  output         io_ipf,
  output         io_isFinish
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
`endif // RANDOMIZE_REG_INIT
  wire [8:0] vpn_vpn0 = io_in_bits_addr[20:12]; // @[EmbeddedTLB.scala 193:54]
  wire [8:0] vpn_vpn1 = io_in_bits_addr[29:21]; // @[EmbeddedTLB.scala 193:54]
  wire [8:0] vpn_vpn2 = io_in_bits_addr[38:30]; // @[EmbeddedTLB.scala 193:54]
  wire [19:0] satp_ppn = io_satp[19:0]; // @[EmbeddedTLB.scala 195:30]
  wire [15:0] satp_asid = io_satp[59:44]; // @[EmbeddedTLB.scala 195:30]
  wire  _T_39 = io_md_0[93:78] == satp_asid; // @[EmbeddedTLB.scala 204:117]
  wire  _T_40 = io_md_0[52] & _T_39; // @[EmbeddedTLB.scala 204:86]
  wire [17:0] _T_57 = {vpn_vpn2,vpn_vpn1}; // @[EmbeddedTLB.scala 204:201]
  wire [26:0] _T_58 = {vpn_vpn2,vpn_vpn1,vpn_vpn0}; // @[EmbeddedTLB.scala 204:201]
  wire [26:0] _T_59 = {9'h1ff,io_md_0[77:60]}; // @[Cat.scala 29:58]
  wire [26:0] _T_60 = _T_59 & io_md_0[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_62 = _T_59 & _T_58; // @[TLB.scala 131:84]
  wire  _T_63 = _T_60 == _T_62; // @[TLB.scala 131:48]
  wire  _T_64 = _T_40 & _T_63; // @[EmbeddedTLB.scala 204:132]
  wire  _T_91 = io_md_1[93:78] == satp_asid; // @[EmbeddedTLB.scala 204:117]
  wire  _T_92 = io_md_1[52] & _T_91; // @[EmbeddedTLB.scala 204:86]
  wire [26:0] _T_111 = {9'h1ff,io_md_1[77:60]}; // @[Cat.scala 29:58]
  wire [26:0] _T_112 = _T_111 & io_md_1[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_114 = _T_111 & _T_58; // @[TLB.scala 131:84]
  wire  _T_115 = _T_112 == _T_114; // @[TLB.scala 131:48]
  wire  _T_116 = _T_92 & _T_115; // @[EmbeddedTLB.scala 204:132]
  wire  _T_143 = io_md_2[93:78] == satp_asid; // @[EmbeddedTLB.scala 204:117]
  wire  _T_144 = io_md_2[52] & _T_143; // @[EmbeddedTLB.scala 204:86]
  wire [26:0] _T_163 = {9'h1ff,io_md_2[77:60]}; // @[Cat.scala 29:58]
  wire [26:0] _T_164 = _T_163 & io_md_2[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_166 = _T_163 & _T_58; // @[TLB.scala 131:84]
  wire  _T_167 = _T_164 == _T_166; // @[TLB.scala 131:48]
  wire  _T_168 = _T_144 & _T_167; // @[EmbeddedTLB.scala 204:132]
  wire  _T_195 = io_md_3[93:78] == satp_asid; // @[EmbeddedTLB.scala 204:117]
  wire  _T_196 = io_md_3[52] & _T_195; // @[EmbeddedTLB.scala 204:86]
  wire [26:0] _T_215 = {9'h1ff,io_md_3[77:60]}; // @[Cat.scala 29:58]
  wire [26:0] _T_216 = _T_215 & io_md_3[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_218 = _T_215 & _T_58; // @[TLB.scala 131:84]
  wire  _T_219 = _T_216 == _T_218; // @[TLB.scala 131:48]
  wire  _T_220 = _T_196 & _T_219; // @[EmbeddedTLB.scala 204:132]
  wire [3:0] hitVec = {_T_220,_T_168,_T_116,_T_64}; // @[EmbeddedTLB.scala 204:211]
  wire  _T_224 = |hitVec; // @[EmbeddedTLB.scala 205:35]
  wire  hit = io_in_valid & _T_224; // @[EmbeddedTLB.scala 205:25]
  wire  _T_226 = ~_T_224; // @[EmbeddedTLB.scala 206:29]
  wire  miss = io_in_valid & _T_226; // @[EmbeddedTLB.scala 206:26]
  reg [63:0] _T_227; // @[LFSR64.scala 25:23]
  wire  _T_230 = _T_227[0] ^ _T_227[1]; // @[LFSR64.scala 26:23]
  wire  _T_232 = _T_230 ^ _T_227[3]; // @[LFSR64.scala 26:33]
  wire  _T_234 = _T_232 ^ _T_227[4]; // @[LFSR64.scala 26:43]
  wire  _T_235 = _T_227 == 64'h0; // @[LFSR64.scala 28:24]
  wire [63:0] _T_237 = {_T_234,_T_227[63:1]}; // @[Cat.scala 29:58]
  wire [3:0] victimWaymask = 4'h1 << _T_227[1:0]; // @[EmbeddedTLB.scala 208:42]
  wire [3:0] waymask = hit ? hitVec : victimWaymask; // @[EmbeddedTLB.scala 209:20]
  wire [120:0] _T_244 = waymask[0] ? io_md_0 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_245 = waymask[1] ? io_md_1 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_246 = waymask[2] ? io_md_2 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_247 = waymask[3] ? io_md_3 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_248 = _T_244 | _T_245; // @[Mux.scala 27:72]
  wire [120:0] _T_249 = _T_248 | _T_246; // @[Mux.scala 27:72]
  wire [120:0] _T_250 = _T_249 | _T_247; // @[Mux.scala 27:72]
  wire [7:0] hitMeta_flag = _T_250[59:52]; // @[EmbeddedTLB.scala 215:70]
  wire [17:0] hitMeta_mask = _T_250[77:60]; // @[EmbeddedTLB.scala 215:70]
  wire [15:0] hitMeta_asid = _T_250[93:78]; // @[EmbeddedTLB.scala 215:70]
  wire [31:0] hitData_pteaddr = _T_250[31:0]; // @[EmbeddedTLB.scala 216:70]
  wire [19:0] hitData_ppn = _T_250[51:32]; // @[EmbeddedTLB.scala 216:70]
  wire  hitFlag_v = hitMeta_flag[0]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_r = hitMeta_flag[1]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_w = hitMeta_flag[2]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_x = hitMeta_flag[3]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_u = hitMeta_flag[4]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_g = hitMeta_flag[5]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_a = hitMeta_flag[6]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_d = hitMeta_flag[7]; // @[EmbeddedTLB.scala 217:38]
  wire  _T_289 = ~hitFlag_a; // @[EmbeddedTLB.scala 221:23]
  wire  _T_294 = hit & _T_289; // @[EmbeddedTLB.scala 221:19]
  wire  _T_314 = io_pf_priviledgeMode == 2'h0; // @[EmbeddedTLB.scala 226:62]
  wire  _T_315 = ~hitFlag_u; // @[EmbeddedTLB.scala 226:75]
  wire  _T_316 = _T_314 & _T_315; // @[EmbeddedTLB.scala 226:72]
  wire  _T_317 = ~_T_316; // @[EmbeddedTLB.scala 226:42]
  wire  _T_318 = hit & _T_317; // @[EmbeddedTLB.scala 226:39]
  wire  _T_319 = io_pf_priviledgeMode == 2'h1; // @[EmbeddedTLB.scala 226:110]
  wire  _T_320 = _T_319 & hitFlag_u; // @[EmbeddedTLB.scala 226:120]
  wire  _T_324 = ~_T_320; // @[EmbeddedTLB.scala 226:90]
  wire  hitCheck = _T_318 & _T_324; // @[EmbeddedTLB.scala 226:87]
  wire  hitExec = hitCheck & hitFlag_x; // @[EmbeddedTLB.scala 227:26]
  wire  _T_329 = ~hitExec; // @[EmbeddedTLB.scala 239:42]
  wire  hitinstrPF = _T_329 & hit; // @[EmbeddedTLB.scala 239:52]
  wire  _T_295 = ~hitinstrPF; // @[EmbeddedTLB.scala 221:69]
  wire  _T_296 = _T_294 & _T_295; // @[EmbeddedTLB.scala 221:66]
  wire  _T_298 = io_pf_loadPF | io_pf_storePF; // @[Bundle.scala 129:23]
  wire  _T_300 = ~_T_298; // @[EmbeddedTLB.scala 221:84]
  wire  hitWB = _T_296 & _T_300; // @[EmbeddedTLB.scala 221:81]
  wire [7:0] _T_310 = {hitFlag_d,hitFlag_a,hitFlag_g,hitFlag_u,hitFlag_x,hitFlag_w,hitFlag_r,hitFlag_v}; // @[EmbeddedTLB.scala 222:79]
  wire [7:0] hitRefillFlag = 8'h40 | _T_310; // @[EmbeddedTLB.scala 222:69]
  wire [39:0] _T_313 = {10'h0,hitData_ppn,2'h0,hitRefillFlag}; // @[Cat.scala 29:58]
  reg [39:0] hitWBStore; // @[Reg.scala 15:16]
  reg [2:0] state; // @[EmbeddedTLB.scala 247:22]
  reg [1:0] level; // @[EmbeddedTLB.scala 248:22]
  reg [63:0] memRespStore; // @[EmbeddedTLB.scala 250:25]
  reg [17:0] missMaskStore; // @[EmbeddedTLB.scala 252:26]
  wire  memRdata_flag_v = io_mem_resp_bits_rdata[0]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_r = io_mem_resp_bits_rdata[1]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_w = io_mem_resp_bits_rdata[2]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_x = io_mem_resp_bits_rdata[3]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_u = io_mem_resp_bits_rdata[4]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_g = io_mem_resp_bits_rdata[5]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_a = io_mem_resp_bits_rdata[6]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_d = io_mem_resp_bits_rdata[7]; // @[EmbeddedTLB.scala 255:49]
  wire [19:0] memRdata_ppn = io_mem_resp_bits_rdata[29:10]; // @[EmbeddedTLB.scala 255:49]
  reg [31:0] raddr; // @[EmbeddedTLB.scala 256:18]
  wire  _T_343 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  reg  alreadyOutFire; // @[Reg.scala 27:20]
  wire  _GEN_2 = _T_343 | alreadyOutFire; // @[Reg.scala 28:19]
  reg  needFlush; // @[EmbeddedTLB.scala 260:26]
  wire  isFlush = needFlush | io_flush; // @[EmbeddedTLB.scala 262:27]
  wire  _T_344 = state != 3'h0; // @[EmbeddedTLB.scala 263:27]
  wire  _T_345 = io_flush & _T_344; // @[EmbeddedTLB.scala 263:17]
  wire  _GEN_3 = _T_345 | needFlush; // @[EmbeddedTLB.scala 263:40]
  wire  _T_347 = _T_343 & needFlush; // @[EmbeddedTLB.scala 264:23]
  wire  _GEN_4 = _T_347 ? 1'h0 : _GEN_3; // @[EmbeddedTLB.scala 264:37]
  reg  missIPF; // @[EmbeddedTLB.scala 266:24]
  wire  _T_348 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_349 = ~io_flush; // @[EmbeddedTLB.scala 271:13]
  wire  _T_350 = _T_349 & hitWB; // @[EmbeddedTLB.scala 271:22]
  wire  _T_352 = miss & _T_349; // @[EmbeddedTLB.scala 275:24]
  wire [31:0] _T_354 = {satp_ppn,vpn_vpn2,3'h0}; // @[Cat.scala 29:58]
  wire  _T_355 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_356 = io_mem_req_ready & io_mem_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_357 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire [7:0] _T_365 = {memRdata_flag_d,memRdata_flag_a,memRdata_flag_g,memRdata_flag_u,memRdata_flag_x,memRdata_flag_w,memRdata_flag_r,memRdata_flag_v}; // @[EmbeddedTLB.scala 292:44]
  wire  _T_375 = io_mem_resp_ready & io_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_376 = _T_365[1] | _T_365[3]; // @[EmbeddedTLB.scala 297:34]
  wire  _T_377 = ~_T_376; // @[EmbeddedTLB.scala 297:21]
  wire  _T_378 = level == 2'h3; // @[EmbeddedTLB.scala 297:58]
  wire  _T_379 = level == 2'h2; // @[EmbeddedTLB.scala 297:73]
  wire  _T_380 = _T_378 | _T_379; // @[EmbeddedTLB.scala 297:65]
  wire  _T_381 = _T_377 & _T_380; // @[EmbeddedTLB.scala 297:49]
  wire  _T_382 = ~_T_365[0]; // @[EmbeddedTLB.scala 298:16]
  wire  _T_383 = ~_T_365[1]; // @[EmbeddedTLB.scala 298:32]
  wire  _T_384 = _T_383 & _T_365[2]; // @[EmbeddedTLB.scala 298:44]
  wire  _T_385 = _T_382 | _T_384; // @[EmbeddedTLB.scala 298:28]
  wire [8:0] _T_417 = _T_378 ? vpn_vpn1 : vpn_vpn0; // @[EmbeddedTLB.scala 311:50]
  wire [31:0] _T_419 = {memRdata_ppn,_T_417,3'h0}; // @[Cat.scala 29:58]
  wire  _GEN_19 = _T_385 | missIPF; // @[EmbeddedTLB.scala 298:60]
  wire  _T_420 = level != 2'h0; // @[EmbeddedTLB.scala 313:27]
  wire  _T_422 = ~_T_365[4]; // @[EmbeddedTLB.scala 314:74]
  wire  _T_423 = _T_314 & _T_422; // @[EmbeddedTLB.scala 314:71]
  wire  _T_424 = ~_T_423; // @[EmbeddedTLB.scala 314:41]
  wire  _T_425 = _T_365[0] & _T_424; // @[EmbeddedTLB.scala 314:38]
  wire  _T_427 = _T_319 & _T_365[4]; // @[EmbeddedTLB.scala 314:120]
  wire  _T_431 = ~_T_427; // @[EmbeddedTLB.scala 314:90]
  wire  _T_432 = _T_425 & _T_431; // @[EmbeddedTLB.scala 314:87]
  wire  _T_433 = _T_432 & _T_365[3]; // @[EmbeddedTLB.scala 315:36]
  wire  _T_438 = ~_T_365[6]; // @[EmbeddedTLB.scala 318:60]
  wire [7:0] _T_456 = {_T_365[7],_T_365[6],_T_365[5],_T_365[4],_T_365[3],_T_365[2],_T_365[1],_T_365[0]}; // @[EmbeddedTLB.scala 320:79]
  wire [7:0] _T_457 = 8'h40 | _T_456; // @[EmbeddedTLB.scala 320:68]
  wire [63:0] _T_458 = io_mem_resp_bits_rdata | 64'h40; // @[EmbeddedTLB.scala 321:50]
  wire  _T_459 = ~_T_433; // @[EmbeddedTLB.scala 323:19]
  wire  _GEN_21 = _T_459 | missIPF; // @[EmbeddedTLB.scala 323:30]
  wire  _GEN_23 = _T_459 ? 1'h0 : 1'h1; // @[EmbeddedTLB.scala 323:30]
  wire  _GEN_28 = _T_420 & _GEN_23; // @[EmbeddedTLB.scala 313:36]
  wire  _GEN_36 = _T_381 ? 1'h0 : _GEN_28; // @[EmbeddedTLB.scala 297:82]
  wire  _GEN_44 = isFlush ? 1'h0 : _GEN_36; // @[EmbeddedTLB.scala 294:24]
  wire [1:0] _T_466 = level - 2'h1; // @[EmbeddedTLB.scala 342:24]
  wire  _GEN_53 = _T_375 & _GEN_44; // @[EmbeddedTLB.scala 293:33]
  wire  _T_467 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_469 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_471 = _T_343 | io_flush; // @[EmbeddedTLB.scala 353:44]
  wire  _T_472 = _T_471 | alreadyOutFire; // @[EmbeddedTLB.scala 353:55]
  wire  _T_473 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_76 = _T_357 & _GEN_53; // @[Conditional.scala 39:67]
  wire  _GEN_87 = _T_355 ? 1'h0 : _GEN_76; // @[Conditional.scala 39:67]
  wire  missMetaRefill = _T_348 ? 1'h0 : _GEN_87; // @[Conditional.scala 40:58]
  wire  cmd = state == 3'h3; // @[EmbeddedTLB.scala 365:23]
  wire  _T_477 = state == 3'h1; // @[EmbeddedTLB.scala 367:31]
  wire  _T_479 = _T_477 | cmd; // @[EmbeddedTLB.scala 367:48]
  wire  _T_480 = ~isFlush; // @[EmbeddedTLB.scala 367:77]
  wire  _T_483 = missMetaRefill & _T_480; // @[EmbeddedTLB.scala 371:50]
  wire  _T_484 = state == 3'h0; // @[EmbeddedTLB.scala 371:82]
  wire  _T_485 = hitWB & _T_484; // @[EmbeddedTLB.scala 371:73]
  wire  _T_487 = _T_485 & _T_480; // @[EmbeddedTLB.scala 371:93]
  wire  _T_488 = _T_483 | _T_487; // @[EmbeddedTLB.scala 371:63]
  reg  _T_489; // @[EmbeddedTLB.scala 371:33]
  reg [3:0] _T_496; // @[EmbeddedTLB.scala 372:60]
  reg [26:0] _T_499; // @[EmbeddedTLB.scala 372:84]
  reg [15:0] _T_501; // @[EmbeddedTLB.scala 373:19]
  reg [17:0] _T_503; // @[EmbeddedTLB.scala 373:72]
  reg [7:0] _T_505; // @[EmbeddedTLB.scala 374:19]
  reg [19:0] _T_507; // @[EmbeddedTLB.scala 374:77]
  reg [31:0] _T_509; // @[EmbeddedTLB.scala 375:22]
  wire [59:0] _T_511 = {_T_505,_T_507,_T_509}; // @[Cat.scala 29:58]
  wire [60:0] _T_513 = {_T_499,_T_501,_T_503}; // @[Cat.scala 29:58]
  wire [31:0] _T_516 = {hitData_ppn,12'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_519 = {2'h3,hitMeta_mask,12'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_520 = _T_516 & _T_519; // @[BitUtils.scala 32:13]
  wire [31:0] _T_521 = ~_T_519; // @[BitUtils.scala 32:38]
  wire [31:0] _T_522 = io_in_bits_addr[31:0] & _T_521; // @[BitUtils.scala 32:36]
  wire [31:0] _T_523 = _T_520 | _T_522; // @[BitUtils.scala 32:25]
  wire [31:0] _T_538 = {memRespStore[29:10],12'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_541 = {2'h3,missMaskStore,12'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_542 = _T_538 & _T_541; // @[BitUtils.scala 32:13]
  wire [31:0] _T_543 = ~_T_541; // @[BitUtils.scala 32:38]
  wire [31:0] _T_544 = io_in_bits_addr[31:0] & _T_543; // @[BitUtils.scala 32:36]
  wire [31:0] _T_545 = _T_542 | _T_544; // @[BitUtils.scala 32:25]
  wire  _T_547 = ~hitWB; // @[EmbeddedTLB.scala 380:45]
  wire  _T_548 = hit & _T_547; // @[EmbeddedTLB.scala 380:42]
  wire  _T_553 = state == 3'h4; // @[EmbeddedTLB.scala 380:97]
  wire  _T_554 = _T_548 ? _T_300 : _T_553; // @[EmbeddedTLB.scala 380:37]
  wire  _T_557 = io_out_ready & _T_484; // @[EmbeddedTLB.scala 382:31]
  wire  _T_558 = ~miss; // @[EmbeddedTLB.scala 382:56]
  wire  _T_559 = _T_557 & _T_558; // @[EmbeddedTLB.scala 382:53]
  wire  _T_561 = _T_559 & _T_547; // @[EmbeddedTLB.scala 382:62]
  wire  _T_562 = _T_561 & io_mdReady; // @[EmbeddedTLB.scala 382:72]
  assign io_in_ready = _T_562 & _T_300; // @[EmbeddedTLB.scala 382:15]
  assign io_out_valid = io_in_valid & _T_554; // @[EmbeddedTLB.scala 380:16]
  assign io_out_bits_addr = hit ? _T_523 : _T_545; // @[EmbeddedTLB.scala 378:15 EmbeddedTLB.scala 379:20]
  assign io_out_bits_user = io_in_bits_user; // @[EmbeddedTLB.scala 378:15]
  assign io_mdWrite_wen = _T_489; // @[TLB.scala 214:14]
  assign io_mdWrite_waymask = _T_496; // @[TLB.scala 216:18]
  assign io_mdWrite_wdata = {_T_513,_T_511}; // @[TLB.scala 217:16]
  assign io_mem_req_valid = _T_479 & _T_480; // @[EmbeddedTLB.scala 367:20]
  assign io_mem_req_bits_addr = hitWB ? hitData_pteaddr : raddr; // @[SimpleBus.scala 64:15]
  assign io_mem_req_bits_cmd = {{3'd0}, cmd}; // @[SimpleBus.scala 65:14]
  assign io_mem_req_bits_wdata = hitWB ? {{24'd0}, hitWBStore} : memRespStore; // @[SimpleBus.scala 67:16]
  assign io_mem_resp_ready = 1'h1; // @[EmbeddedTLB.scala 368:21]
  assign io_pf_loadPF = 1'h0; // @[EmbeddedTLB.scala 199:13 EmbeddedTLB.scala 236:16]
  assign io_pf_storePF = 1'h0; // @[EmbeddedTLB.scala 200:14 EmbeddedTLB.scala 237:17]
  assign io_ipf = hit ? hitinstrPF : missIPF; // @[EmbeddedTLB.scala 384:10]
  assign io_isFinish = _T_343 | _T_298; // @[EmbeddedTLB.scala 385:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _T_227 = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  hitWBStore = _RAND_1[39:0];
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  level = _RAND_3[1:0];
  _RAND_4 = {2{`RANDOM}};
  memRespStore = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  missMaskStore = _RAND_5[17:0];
  _RAND_6 = {1{`RANDOM}};
  raddr = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  alreadyOutFire = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  needFlush = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  missIPF = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _T_489 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_496 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  _T_499 = _RAND_12[26:0];
  _RAND_13 = {1{`RANDOM}};
  _T_501 = _RAND_13[15:0];
  _RAND_14 = {1{`RANDOM}};
  _T_503 = _RAND_14[17:0];
  _RAND_15 = {1{`RANDOM}};
  _T_505 = _RAND_15[7:0];
  _RAND_16 = {1{`RANDOM}};
  _T_507 = _RAND_16[19:0];
  _RAND_17 = {1{`RANDOM}};
  _T_509 = _RAND_17[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_227 <= 64'h1234567887654321;
    end else if (_T_235) begin
      _T_227 <= 64'h1;
    end else begin
      _T_227 <= _T_237;
    end
    if (hitWB) begin
      hitWBStore <= _T_313;
    end
    if (reset) begin
      state <= 3'h0;
    end else if (_T_348) begin
      if (_T_350) begin
        state <= 3'h3;
      end else if (_T_352) begin
        state <= 3'h1;
      end
    end else if (_T_355) begin
      if (isFlush) begin
        state <= 3'h0;
      end else if (_T_356) begin
        state <= 3'h2;
      end
    end else if (_T_357) begin
      if (_T_375) begin
        if (isFlush) begin
          state <= 3'h0;
        end else if (_T_381) begin
          if (_T_385) begin
            state <= 3'h4;
          end else begin
            state <= 3'h1;
          end
        end else if (_T_420) begin
          if (_T_459) begin
            state <= 3'h4;
          end else if (_T_438) begin
            state <= 3'h3;
          end else begin
            state <= 3'h4;
          end
        end
      end
    end else if (_T_467) begin
      if (isFlush) begin
        state <= 3'h0;
      end else if (_T_356) begin
        state <= 3'h4;
      end
    end else if (_T_469) begin
      if (_T_472) begin
        state <= 3'h0;
      end
    end else if (_T_473) begin
      state <= 3'h0;
    end
    if (reset) begin
      level <= 2'h3;
    end else if (_T_348) begin
      if (!(_T_350)) begin
        if (_T_352) begin
          level <= 2'h3;
        end
      end
    end else if (!(_T_355)) begin
      if (_T_357) begin
        if (_T_375) begin
          level <= _T_466;
        end
      end
    end
    if (!(_T_348)) begin
      if (!(_T_355)) begin
        if (_T_357) begin
          if (_T_375) begin
            if (!(isFlush)) begin
              if (!(_T_381)) begin
                if (_T_420) begin
                  memRespStore <= _T_458;
                end
              end
            end
          end
        end
      end
    end
    if (!(_T_348)) begin
      if (!(_T_355)) begin
        if (_T_357) begin
          if (_T_375) begin
            if (!(isFlush)) begin
              if (!(_T_381)) begin
                if (_T_420) begin
                  if (_T_348) begin
                    missMaskStore <= 18'h3ffff;
                  end else if (_T_355) begin
                    missMaskStore <= 18'h3ffff;
                  end else if (_T_357) begin
                    if (_T_375) begin
                      if (isFlush) begin
                        missMaskStore <= 18'h3ffff;
                      end else if (_T_381) begin
                        missMaskStore <= 18'h3ffff;
                      end else if (_T_420) begin
                        if (_T_378) begin
                          missMaskStore <= 18'h0;
                        end else if (_T_379) begin
                          missMaskStore <= 18'h3fe00;
                        end else begin
                          missMaskStore <= 18'h3ffff;
                        end
                      end else begin
                        missMaskStore <= 18'h3ffff;
                      end
                    end else begin
                      missMaskStore <= 18'h3ffff;
                    end
                  end else begin
                    missMaskStore <= 18'h3ffff;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_348) begin
      if (!(_T_350)) begin
        if (_T_352) begin
          raddr <= _T_354;
        end
      end
    end else if (!(_T_355)) begin
      if (_T_357) begin
        if (_T_375) begin
          if (!(isFlush)) begin
            if (_T_381) begin
              if (!(_T_385)) begin
                raddr <= _T_419;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      alreadyOutFire <= 1'h0;
    end else if (_T_348) begin
      if (_T_350) begin
        alreadyOutFire <= 1'h0;
      end else if (_T_352) begin
        alreadyOutFire <= 1'h0;
      end else begin
        alreadyOutFire <= _GEN_2;
      end
    end else if (_T_355) begin
      alreadyOutFire <= _GEN_2;
    end else if (_T_357) begin
      alreadyOutFire <= _GEN_2;
    end else if (_T_467) begin
      alreadyOutFire <= _GEN_2;
    end else if (_T_469) begin
      if (_T_472) begin
        alreadyOutFire <= 1'h0;
      end else begin
        alreadyOutFire <= _GEN_2;
      end
    end else begin
      alreadyOutFire <= _GEN_2;
    end
    if (reset) begin
      needFlush <= 1'h0;
    end else if (_T_348) begin
      if (_T_350) begin
        needFlush <= 1'h0;
      end else if (_T_352) begin
        needFlush <= 1'h0;
      end else if (_T_347) begin
        needFlush <= 1'h0;
      end else begin
        needFlush <= _GEN_3;
      end
    end else if (_T_355) begin
      if (isFlush) begin
        needFlush <= 1'h0;
      end else if (_T_347) begin
        needFlush <= 1'h0;
      end else begin
        needFlush <= _GEN_3;
      end
    end else if (_T_357) begin
      if (_T_375) begin
        if (isFlush) begin
          needFlush <= 1'h0;
        end else if (_T_347) begin
          needFlush <= 1'h0;
        end else begin
          needFlush <= _GEN_3;
        end
      end else if (_T_347) begin
        needFlush <= 1'h0;
      end else begin
        needFlush <= _GEN_3;
      end
    end else if (_T_467) begin
      if (isFlush) begin
        needFlush <= 1'h0;
      end else begin
        needFlush <= _GEN_4;
      end
    end else begin
      needFlush <= _GEN_4;
    end
    if (reset) begin
      missIPF <= 1'h0;
    end else if (!(_T_348)) begin
      if (!(_T_355)) begin
        if (_T_357) begin
          if (_T_375) begin
            if (!(isFlush)) begin
              if (_T_381) begin
                missIPF <= _GEN_19;
              end else if (_T_420) begin
                missIPF <= _GEN_21;
              end
            end
          end
        end else if (!(_T_467)) begin
          if (_T_469) begin
            if (_T_472) begin
              missIPF <= 1'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      _T_489 <= 1'h0;
    end else begin
      _T_489 <= _T_488;
    end
    if (hit) begin
      _T_496 <= hitVec;
    end else begin
      _T_496 <= victimWaymask;
    end
    _T_499 <= {_T_57,vpn_vpn0};
    if (hitWB) begin
      _T_501 <= hitMeta_asid;
    end else begin
      _T_501 <= satp_asid;
    end
    if (hitWB) begin
      _T_503 <= hitMeta_mask;
    end else if (_T_348) begin
      _T_503 <= 18'h3ffff;
    end else if (_T_355) begin
      _T_503 <= 18'h3ffff;
    end else if (_T_357) begin
      if (_T_375) begin
        if (isFlush) begin
          _T_503 <= 18'h3ffff;
        end else if (_T_381) begin
          _T_503 <= 18'h3ffff;
        end else if (_T_420) begin
          if (_T_378) begin
            _T_503 <= 18'h0;
          end else if (_T_379) begin
            _T_503 <= 18'h3fe00;
          end else begin
            _T_503 <= 18'h3ffff;
          end
        end else begin
          _T_503 <= 18'h3ffff;
        end
      end else begin
        _T_503 <= 18'h3ffff;
      end
    end else begin
      _T_503 <= 18'h3ffff;
    end
    if (hitWB) begin
      _T_505 <= hitRefillFlag;
    end else if (_T_348) begin
      _T_505 <= 8'h0;
    end else if (_T_355) begin
      _T_505 <= 8'h0;
    end else if (_T_357) begin
      if (_T_375) begin
        if (isFlush) begin
          _T_505 <= 8'h0;
        end else if (_T_381) begin
          _T_505 <= 8'h0;
        end else if (_T_420) begin
          _T_505 <= _T_457;
        end else begin
          _T_505 <= 8'h0;
        end
      end else begin
        _T_505 <= 8'h0;
      end
    end else begin
      _T_505 <= 8'h0;
    end
    if (hitWB) begin
      _T_507 <= hitData_ppn;
    end else begin
      _T_507 <= memRdata_ppn;
    end
    if (hitWB) begin
      _T_509 <= hitData_pteaddr;
    end else begin
      _T_509 <= raddr;
    end
  end
endmodule
module EmbeddedTLBMD(
  input          clock,
  input          reset,
  output [120:0] io_tlbmd_0,
  output [120:0] io_tlbmd_1,
  output [120:0] io_tlbmd_2,
  output [120:0] io_tlbmd_3,
  input          io_write_wen,
  input  [3:0]   io_write_waymask,
  input  [120:0] io_write_wdata,
  output         io_ready
);
`ifdef RANDOMIZE_MEM_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  reg [120:0] tlbmd_0 [0:0]; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_0__T_data; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_0__T_addr; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_0__T_6_data; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_0__T_6_addr; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_0__T_6_mask; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_0__T_6_en; // @[EmbeddedTLB.scala 38:18]
  reg [120:0] tlbmd_1 [0:0]; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_1__T_data; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_1__T_addr; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_1__T_6_data; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_1__T_6_addr; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_1__T_6_mask; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_1__T_6_en; // @[EmbeddedTLB.scala 38:18]
  reg [120:0] tlbmd_2 [0:0]; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_2__T_data; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_2__T_addr; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_2__T_6_data; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_2__T_6_addr; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_2__T_6_mask; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_2__T_6_en; // @[EmbeddedTLB.scala 38:18]
  reg [120:0] tlbmd_3 [0:0]; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_3__T_data; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_3__T_addr; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_3__T_6_data; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_3__T_6_addr; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_3__T_6_mask; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_3__T_6_en; // @[EmbeddedTLB.scala 38:18]
  reg  resetState; // @[EmbeddedTLB.scala 42:27]
  wire  _GEN_1 = resetState ? 1'h0 : resetState; // @[EmbeddedTLB.scala 44:22]
  wire [3:0] waymask = resetState ? 4'hf : io_write_waymask; // @[EmbeddedTLB.scala 53:20]
  assign tlbmd_0__T_addr = 1'h0;
  assign tlbmd_0__T_data = tlbmd_0[tlbmd_0__T_addr]; // @[EmbeddedTLB.scala 38:18]
  assign tlbmd_0__T_6_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_0__T_6_addr = 1'h0;
  assign tlbmd_0__T_6_mask = waymask[0];
  assign tlbmd_0__T_6_en = resetState | io_write_wen;
  assign tlbmd_1__T_addr = 1'h0;
  assign tlbmd_1__T_data = tlbmd_1[tlbmd_1__T_addr]; // @[EmbeddedTLB.scala 38:18]
  assign tlbmd_1__T_6_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_1__T_6_addr = 1'h0;
  assign tlbmd_1__T_6_mask = waymask[1];
  assign tlbmd_1__T_6_en = resetState | io_write_wen;
  assign tlbmd_2__T_addr = 1'h0;
  assign tlbmd_2__T_data = tlbmd_2[tlbmd_2__T_addr]; // @[EmbeddedTLB.scala 38:18]
  assign tlbmd_2__T_6_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_2__T_6_addr = 1'h0;
  assign tlbmd_2__T_6_mask = waymask[2];
  assign tlbmd_2__T_6_en = resetState | io_write_wen;
  assign tlbmd_3__T_addr = 1'h0;
  assign tlbmd_3__T_data = tlbmd_3[tlbmd_3__T_addr]; // @[EmbeddedTLB.scala 38:18]
  assign tlbmd_3__T_6_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_3__T_6_addr = 1'h0;
  assign tlbmd_3__T_6_mask = waymask[3];
  assign tlbmd_3__T_6_en = resetState | io_write_wen;
  assign io_tlbmd_0 = tlbmd_0__T_data; // @[EmbeddedTLB.scala 39:12]
  assign io_tlbmd_1 = tlbmd_1__T_data; // @[EmbeddedTLB.scala 39:12]
  assign io_tlbmd_2 = tlbmd_2__T_data; // @[EmbeddedTLB.scala 39:12]
  assign io_tlbmd_3 = tlbmd_3__T_data; // @[EmbeddedTLB.scala 39:12]
  assign io_ready = ~resetState; // @[EmbeddedTLB.scala 59:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {4{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_0[initvar] = _RAND_0[120:0];
  _RAND_1 = {4{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_1[initvar] = _RAND_1[120:0];
  _RAND_2 = {4{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_2[initvar] = _RAND_2[120:0];
  _RAND_3 = {4{`RANDOM}};
  for (initvar = 0; initvar < 1; initvar = initvar+1)
    tlbmd_3[initvar] = _RAND_3[120:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  resetState = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(tlbmd_0__T_6_en & tlbmd_0__T_6_mask) begin
      tlbmd_0[tlbmd_0__T_6_addr] <= tlbmd_0__T_6_data; // @[EmbeddedTLB.scala 38:18]
    end
    if(tlbmd_1__T_6_en & tlbmd_1__T_6_mask) begin
      tlbmd_1[tlbmd_1__T_6_addr] <= tlbmd_1__T_6_data; // @[EmbeddedTLB.scala 38:18]
    end
    if(tlbmd_2__T_6_en & tlbmd_2__T_6_mask) begin
      tlbmd_2[tlbmd_2__T_6_addr] <= tlbmd_2__T_6_data; // @[EmbeddedTLB.scala 38:18]
    end
    if(tlbmd_3__T_6_en & tlbmd_3__T_6_mask) begin
      tlbmd_3[tlbmd_3__T_6_addr] <= tlbmd_3__T_6_data; // @[EmbeddedTLB.scala 38:18]
    end
    resetState <= reset | _GEN_1;
  end
endmodule
module EmbeddedTLB(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [38:0] io_in_req_bits_addr,
  input  [86:0] io_in_req_bits_user,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  output [86:0] io_in_resp_bits_user,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [86:0] io_out_req_bits_user,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [63:0] io_out_resp_bits_rdata,
  input  [86:0] io_out_resp_bits_user,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [31:0] io_mem_req_bits_addr,
  output [3:0]  io_mem_req_bits_cmd,
  output [63:0] io_mem_req_bits_wdata,
  input         io_mem_resp_valid,
  input  [63:0] io_mem_resp_bits_rdata,
  input         io_flush,
  input  [1:0]  io_csrMMU_priviledgeMode,
  input         io_cacheEmpty,
  output        io_ipf,
  input  [63:0] CSRSATP,
  input         MOUFlushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [95:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  tlbExec_clock; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_reset; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_in_ready; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_in_valid; // @[EmbeddedTLB.scala 80:23]
  wire [38:0] tlbExec_io_in_bits_addr; // @[EmbeddedTLB.scala 80:23]
  wire [86:0] tlbExec_io_in_bits_user; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_out_ready; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_out_valid; // @[EmbeddedTLB.scala 80:23]
  wire [31:0] tlbExec_io_out_bits_addr; // @[EmbeddedTLB.scala 80:23]
  wire [86:0] tlbExec_io_out_bits_user; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_md_0; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_md_1; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_md_2; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_md_3; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mdWrite_wen; // @[EmbeddedTLB.scala 80:23]
  wire [3:0] tlbExec_io_mdWrite_waymask; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_mdWrite_wdata; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mdReady; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mem_req_ready; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mem_req_valid; // @[EmbeddedTLB.scala 80:23]
  wire [31:0] tlbExec_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 80:23]
  wire [3:0] tlbExec_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 80:23]
  wire [63:0] tlbExec_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mem_resp_ready; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mem_resp_valid; // @[EmbeddedTLB.scala 80:23]
  wire [63:0] tlbExec_io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_flush; // @[EmbeddedTLB.scala 80:23]
  wire [63:0] tlbExec_io_satp; // @[EmbeddedTLB.scala 80:23]
  wire [1:0] tlbExec_io_pf_priviledgeMode; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_pf_loadPF; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_pf_storePF; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_ipf; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_isFinish; // @[EmbeddedTLB.scala 80:23]
  wire  mdTLB_clock; // @[EmbeddedTLB.scala 82:21]
  wire  mdTLB_reset; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_tlbmd_0; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_tlbmd_1; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_tlbmd_2; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_tlbmd_3; // @[EmbeddedTLB.scala 82:21]
  wire  mdTLB_io_write_wen; // @[EmbeddedTLB.scala 82:21]
  wire [3:0] mdTLB_io_write_waymask; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_write_wdata; // @[EmbeddedTLB.scala 82:21]
  wire  mdTLB_io_ready; // @[EmbeddedTLB.scala 82:21]
  reg [120:0] _T__0; // @[Reg.scala 15:16]
  reg [120:0] _T__1; // @[Reg.scala 15:16]
  reg [120:0] _T__2; // @[Reg.scala 15:16]
  reg [120:0] _T__3; // @[Reg.scala 15:16]
  wire  mdUpdate = io_in_req_valid & tlbExec_io_in_ready; // @[EmbeddedTLB.scala 114:26]
  wire  _T_14 = CSRSATP[63:60] == 4'h8; // @[EmbeddedTLB.scala 102:49]
  wire  _T_15 = io_csrMMU_priviledgeMode < 2'h3; // @[EmbeddedTLB.scala 102:86]
  wire  vmEnable = _T_14 & _T_15; // @[EmbeddedTLB.scala 102:57]
  reg  _T_16; // @[EmbeddedTLB.scala 105:24]
  wire  _GEN_4 = tlbExec_io_isFinish ? 1'h0 : _T_16; // @[EmbeddedTLB.scala 106:25]
  wire  _T_18 = mdUpdate & vmEnable; // @[EmbeddedTLB.scala 107:37]
  wire  _GEN_5 = _T_18 | _GEN_4; // @[EmbeddedTLB.scala 107:50]
  reg [38:0] _T_20_addr; // @[Reg.scala 15:16]
  reg [86:0] _T_20_user; // @[Reg.scala 15:16]
  wire  _T_22 = ~vmEnable; // @[EmbeddedTLB.scala 123:8]
  wire  _GEN_13 = _T_22 | io_out_req_ready; // @[EmbeddedTLB.scala 123:19]
  wire  _GEN_14 = _T_22 ? io_in_req_valid : tlbExec_io_out_valid; // @[EmbeddedTLB.scala 123:19]
  wire  _T_24 = tlbExec_io_ipf & vmEnable; // @[EmbeddedTLB.scala 152:26]
  wire  _T_25 = io_cacheEmpty & io_in_resp_ready; // @[EmbeddedTLB.scala 153:45]
  wire  _T_27 = _T_24 & io_cacheEmpty; // @[EmbeddedTLB.scala 157:38]
  EmbeddedTLBExec tlbExec ( // @[EmbeddedTLB.scala 80:23]
    .clock(tlbExec_clock),
    .reset(tlbExec_reset),
    .io_in_ready(tlbExec_io_in_ready),
    .io_in_valid(tlbExec_io_in_valid),
    .io_in_bits_addr(tlbExec_io_in_bits_addr),
    .io_in_bits_user(tlbExec_io_in_bits_user),
    .io_out_ready(tlbExec_io_out_ready),
    .io_out_valid(tlbExec_io_out_valid),
    .io_out_bits_addr(tlbExec_io_out_bits_addr),
    .io_out_bits_user(tlbExec_io_out_bits_user),
    .io_md_0(tlbExec_io_md_0),
    .io_md_1(tlbExec_io_md_1),
    .io_md_2(tlbExec_io_md_2),
    .io_md_3(tlbExec_io_md_3),
    .io_mdWrite_wen(tlbExec_io_mdWrite_wen),
    .io_mdWrite_waymask(tlbExec_io_mdWrite_waymask),
    .io_mdWrite_wdata(tlbExec_io_mdWrite_wdata),
    .io_mdReady(tlbExec_io_mdReady),
    .io_mem_req_ready(tlbExec_io_mem_req_ready),
    .io_mem_req_valid(tlbExec_io_mem_req_valid),
    .io_mem_req_bits_addr(tlbExec_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(tlbExec_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(tlbExec_io_mem_req_bits_wdata),
    .io_mem_resp_ready(tlbExec_io_mem_resp_ready),
    .io_mem_resp_valid(tlbExec_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(tlbExec_io_mem_resp_bits_rdata),
    .io_flush(tlbExec_io_flush),
    .io_satp(tlbExec_io_satp),
    .io_pf_priviledgeMode(tlbExec_io_pf_priviledgeMode),
    .io_pf_loadPF(tlbExec_io_pf_loadPF),
    .io_pf_storePF(tlbExec_io_pf_storePF),
    .io_ipf(tlbExec_io_ipf),
    .io_isFinish(tlbExec_io_isFinish)
  );
  EmbeddedTLBMD mdTLB ( // @[EmbeddedTLB.scala 82:21]
    .clock(mdTLB_clock),
    .reset(mdTLB_reset),
    .io_tlbmd_0(mdTLB_io_tlbmd_0),
    .io_tlbmd_1(mdTLB_io_tlbmd_1),
    .io_tlbmd_2(mdTLB_io_tlbmd_2),
    .io_tlbmd_3(mdTLB_io_tlbmd_3),
    .io_write_wen(mdTLB_io_write_wen),
    .io_write_waymask(mdTLB_io_write_waymask),
    .io_write_wdata(mdTLB_io_write_wdata),
    .io_ready(mdTLB_io_ready)
  );
  assign io_in_req_ready = _T_22 ? io_out_req_ready : tlbExec_io_in_ready; // @[EmbeddedTLB.scala 110:16 EmbeddedTLB.scala 127:21]
  assign io_in_resp_valid = _T_27 | io_out_resp_valid; // @[EmbeddedTLB.scala 138:15 EmbeddedTLB.scala 158:24]
  assign io_in_resp_bits_rdata = _T_27 ? 64'h0 : io_out_resp_bits_rdata; // @[EmbeddedTLB.scala 138:15 EmbeddedTLB.scala 159:29]
  assign io_in_resp_bits_user = _T_27 ? tlbExec_io_in_bits_user : io_out_resp_bits_user; // @[EmbeddedTLB.scala 138:15 EmbeddedTLB.scala 161:34]
  assign io_out_req_valid = _T_24 ? 1'h0 : _GEN_14; // @[EmbeddedTLB.scala 126:22 EmbeddedTLB.scala 136:23 EmbeddedTLB.scala 154:24]
  assign io_out_req_bits_addr = _T_22 ? io_in_req_bits_addr[31:0] : tlbExec_io_out_bits_addr; // @[EmbeddedTLB.scala 128:26 EmbeddedTLB.scala 136:23]
  assign io_out_req_bits_user = _T_22 ? io_in_req_bits_user : tlbExec_io_out_bits_user; // @[EmbeddedTLB.scala 133:32 EmbeddedTLB.scala 136:23]
  assign io_out_resp_ready = io_in_resp_ready; // @[EmbeddedTLB.scala 138:15]
  assign io_mem_req_valid = tlbExec_io_mem_req_valid; // @[EmbeddedTLB.scala 87:18]
  assign io_mem_req_bits_addr = tlbExec_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 87:18]
  assign io_mem_req_bits_cmd = tlbExec_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 87:18]
  assign io_mem_req_bits_wdata = tlbExec_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 87:18]
  assign io_ipf = _T_27 & tlbExec_io_ipf; // @[EmbeddedTLB.scala 94:10 EmbeddedTLB.scala 162:14]
  assign tlbExec_clock = clock;
  assign tlbExec_reset = reset;
  assign tlbExec_io_in_valid = _T_16; // @[EmbeddedTLB.scala 112:17]
  assign tlbExec_io_in_bits_addr = _T_20_addr; // @[EmbeddedTLB.scala 111:16]
  assign tlbExec_io_in_bits_user = _T_20_user; // @[EmbeddedTLB.scala 111:16]
  assign tlbExec_io_out_ready = _T_24 ? _T_25 : _GEN_13; // @[EmbeddedTLB.scala 124:26 EmbeddedTLB.scala 136:23 EmbeddedTLB.scala 153:28]
  assign tlbExec_io_md_0 = _T__0; // @[EmbeddedTLB.scala 89:17]
  assign tlbExec_io_md_1 = _T__1; // @[EmbeddedTLB.scala 89:17]
  assign tlbExec_io_md_2 = _T__2; // @[EmbeddedTLB.scala 89:17]
  assign tlbExec_io_md_3 = _T__3; // @[EmbeddedTLB.scala 89:17]
  assign tlbExec_io_mdReady = mdTLB_io_ready; // @[EmbeddedTLB.scala 90:22]
  assign tlbExec_io_mem_req_ready = io_mem_req_ready; // @[EmbeddedTLB.scala 87:18]
  assign tlbExec_io_mem_resp_valid = io_mem_resp_valid; // @[EmbeddedTLB.scala 87:18]
  assign tlbExec_io_mem_resp_bits_rdata = io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 87:18]
  assign tlbExec_io_flush = io_flush; // @[EmbeddedTLB.scala 85:20]
  assign tlbExec_io_satp = CSRSATP; // @[EmbeddedTLB.scala 86:19]
  assign tlbExec_io_pf_priviledgeMode = io_csrMMU_priviledgeMode; // @[EmbeddedTLB.scala 88:17]
  assign mdTLB_clock = clock;
  assign mdTLB_reset = reset | MOUFlushTLB; // @[EmbeddedTLB.scala 99:15]
  assign mdTLB_io_write_wen = tlbExec_io_mdWrite_wen; // @[EmbeddedTLB.scala 92:18]
  assign mdTLB_io_write_waymask = tlbExec_io_mdWrite_waymask; // @[EmbeddedTLB.scala 92:18]
  assign mdTLB_io_write_wdata = tlbExec_io_mdWrite_wdata; // @[EmbeddedTLB.scala 92:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  _T__0 = _RAND_0[120:0];
  _RAND_1 = {4{`RANDOM}};
  _T__1 = _RAND_1[120:0];
  _RAND_2 = {4{`RANDOM}};
  _T__2 = _RAND_2[120:0];
  _RAND_3 = {4{`RANDOM}};
  _T__3 = _RAND_3[120:0];
  _RAND_4 = {1{`RANDOM}};
  _T_16 = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  _T_20_addr = _RAND_5[38:0];
  _RAND_6 = {3{`RANDOM}};
  _T_20_user = _RAND_6[86:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (mdUpdate) begin
      _T__0 <= mdTLB_io_tlbmd_0;
    end
    if (mdUpdate) begin
      _T__1 <= mdTLB_io_tlbmd_1;
    end
    if (mdUpdate) begin
      _T__2 <= mdTLB_io_tlbmd_2;
    end
    if (mdUpdate) begin
      _T__3 <= mdTLB_io_tlbmd_3;
    end
    if (reset) begin
      _T_16 <= 1'h0;
    end else if (io_flush) begin
      _T_16 <= 1'h0;
    end else begin
      _T_16 <= _GEN_5;
    end
    if (mdUpdate) begin
      _T_20_addr <= io_in_req_bits_addr;
    end
    if (mdUpdate) begin
      _T_20_user <= io_in_req_bits_user;
    end
  end
endmodule
module CacheStage1(
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [86:0] io_in_bits_user,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [86:0] io_out_bits_req_user,
  input         io_metaReadBus_req_ready,
  output        io_metaReadBus_req_valid,
  output [6:0]  io_metaReadBus_req_bits_setIdx,
  input  [18:0] io_metaReadBus_resp_data_0_tag,
  input         io_metaReadBus_resp_data_0_valid,
  input         io_metaReadBus_resp_data_0_dirty,
  input  [18:0] io_metaReadBus_resp_data_1_tag,
  input         io_metaReadBus_resp_data_1_valid,
  input         io_metaReadBus_resp_data_1_dirty,
  input  [18:0] io_metaReadBus_resp_data_2_tag,
  input         io_metaReadBus_resp_data_2_valid,
  input         io_metaReadBus_resp_data_2_dirty,
  input  [18:0] io_metaReadBus_resp_data_3_tag,
  input         io_metaReadBus_resp_data_3_valid,
  input         io_metaReadBus_resp_data_3_dirty,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [9:0]  io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data
);
  wire  _T_35 = io_in_valid & io_metaReadBus_req_ready; // @[Cache.scala 133:31]
  wire  _T_37 = ~io_in_valid; // @[Cache.scala 134:19]
  wire  _T_38 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_39 = _T_37 | _T_38; // @[Cache.scala 134:32]
  wire  _T_40 = _T_39 & io_metaReadBus_req_ready; // @[Cache.scala 134:50]
  assign io_in_ready = _T_40 & io_dataReadBus_req_ready; // @[Cache.scala 134:15]
  assign io_out_valid = _T_35 & io_dataReadBus_req_ready; // @[Cache.scala 133:16]
  assign io_out_bits_req_addr = io_in_bits_addr; // @[Cache.scala 132:19]
  assign io_out_bits_req_user = io_in_bits_user; // @[Cache.scala 132:19]
  assign io_metaReadBus_req_valid = io_in_valid & io_out_ready; // @[SRAMTemplate.scala 53:20]
  assign io_metaReadBus_req_bits_setIdx = io_in_bits_addr[12:6]; // @[SRAMTemplate.scala 26:17]
  assign io_dataReadBus_req_valid = io_in_valid & io_out_ready; // @[SRAMTemplate.scala 53:20]
  assign io_dataReadBus_req_bits_setIdx = {io_in_bits_addr[12:6],io_in_bits_addr[5:3]}; // @[SRAMTemplate.scala 26:17]
endmodule
module CacheStage2(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [86:0] io_in_bits_req_user,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [86:0] io_out_bits_req_user,
  output [18:0] io_out_bits_metas_0_tag,
  output        io_out_bits_metas_0_valid,
  output        io_out_bits_metas_0_dirty,
  output [18:0] io_out_bits_metas_1_tag,
  output        io_out_bits_metas_1_valid,
  output        io_out_bits_metas_1_dirty,
  output [18:0] io_out_bits_metas_2_tag,
  output        io_out_bits_metas_2_valid,
  output        io_out_bits_metas_2_dirty,
  output [18:0] io_out_bits_metas_3_tag,
  output        io_out_bits_metas_3_valid,
  output        io_out_bits_metas_3_dirty,
  output [63:0] io_out_bits_datas_0_data,
  output [63:0] io_out_bits_datas_1_data,
  output [63:0] io_out_bits_datas_2_data,
  output [63:0] io_out_bits_datas_3_data,
  output        io_out_bits_hit,
  output [3:0]  io_out_bits_waymask,
  output        io_out_bits_mmio,
  output        io_out_bits_isForwardData,
  output [63:0] io_out_bits_forwardData_data_data,
  output [3:0]  io_out_bits_forwardData_waymask,
  input  [18:0] io_metaReadResp_0_tag,
  input         io_metaReadResp_0_valid,
  input         io_metaReadResp_0_dirty,
  input  [18:0] io_metaReadResp_1_tag,
  input         io_metaReadResp_1_valid,
  input         io_metaReadResp_1_dirty,
  input  [18:0] io_metaReadResp_2_tag,
  input         io_metaReadResp_2_valid,
  input         io_metaReadResp_2_dirty,
  input  [18:0] io_metaReadResp_3_tag,
  input         io_metaReadResp_3_valid,
  input         io_metaReadResp_3_dirty,
  input  [63:0] io_dataReadResp_0_data,
  input  [63:0] io_dataReadResp_1_data,
  input  [63:0] io_dataReadResp_2_data,
  input  [63:0] io_dataReadResp_3_data,
  input         io_metaWriteBus_req_valid,
  input  [6:0]  io_metaWriteBus_req_bits_setIdx,
  input  [18:0] io_metaWriteBus_req_bits_data_tag,
  input         io_metaWriteBus_req_bits_data_dirty,
  input  [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_dataWriteBus_req_valid,
  input  [9:0]  io_dataWriteBus_req_bits_setIdx,
  input  [63:0] io_dataWriteBus_req_bits_data_data,
  input  [3:0]  io_dataWriteBus_req_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 162:31]
  wire [6:0] addr_index = io_in_bits_req_addr[12:6]; // @[Cache.scala 162:31]
  wire [18:0] addr_tag = io_in_bits_req_addr[31:13]; // @[Cache.scala 162:31]
  wire  _T_5 = io_in_valid & io_metaWriteBus_req_valid; // @[Cache.scala 164:35]
  wire  _T_12 = io_metaWriteBus_req_bits_setIdx == addr_index; // @[Cache.scala 164:99]
  wire  isForwardMeta = _T_5 & _T_12; // @[Cache.scala 164:64]
  reg  isForwardMetaReg; // @[Cache.scala 165:33]
  wire  _GEN_0 = isForwardMeta | isForwardMetaReg; // @[Cache.scala 166:24]
  wire  _T_13 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire  _T_14 = ~io_in_valid; // @[Cache.scala 167:25]
  wire  _T_15 = _T_13 | _T_14; // @[Cache.scala 167:22]
  reg [18:0] forwardMetaReg_data_tag; // @[Reg.scala 15:16]
  reg  forwardMetaReg_data_dirty; // @[Reg.scala 15:16]
  reg [3:0] forwardMetaReg_waymask; // @[Reg.scala 15:16]
  wire [3:0] _GEN_2 = isForwardMeta ? io_metaWriteBus_req_bits_waymask : forwardMetaReg_waymask; // @[Reg.scala 16:19]
  wire  _GEN_3 = isForwardMeta ? io_metaWriteBus_req_bits_data_dirty : forwardMetaReg_data_dirty; // @[Reg.scala 16:19]
  wire [18:0] _GEN_5 = isForwardMeta ? io_metaWriteBus_req_bits_data_tag : forwardMetaReg_data_tag; // @[Reg.scala 16:19]
  wire  pickForwardMeta = isForwardMetaReg | isForwardMeta; // @[Cache.scala 171:42]
  wire  forwardWaymask_0 = _GEN_2[0]; // @[Cache.scala 173:61]
  wire  forwardWaymask_1 = _GEN_2[1]; // @[Cache.scala 173:61]
  wire  forwardWaymask_2 = _GEN_2[2]; // @[Cache.scala 173:61]
  wire  forwardWaymask_3 = _GEN_2[3]; // @[Cache.scala 173:61]
  wire  _T_16 = pickForwardMeta & forwardWaymask_0; // @[Cache.scala 175:39]
  wire [18:0] metaWay_0_tag = _T_16 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 175:22]
  wire  metaWay_0_valid = _T_16 | io_metaReadResp_0_valid; // @[Cache.scala 175:22]
  wire  _T_18 = pickForwardMeta & forwardWaymask_1; // @[Cache.scala 175:39]
  wire [18:0] metaWay_1_tag = _T_18 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 175:22]
  wire  metaWay_1_valid = _T_18 | io_metaReadResp_1_valid; // @[Cache.scala 175:22]
  wire  _T_20 = pickForwardMeta & forwardWaymask_2; // @[Cache.scala 175:39]
  wire [18:0] metaWay_2_tag = _T_20 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 175:22]
  wire  metaWay_2_valid = _T_20 | io_metaReadResp_2_valid; // @[Cache.scala 175:22]
  wire  _T_22 = pickForwardMeta & forwardWaymask_3; // @[Cache.scala 175:39]
  wire [18:0] metaWay_3_tag = _T_22 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 175:22]
  wire  metaWay_3_valid = _T_22 | io_metaReadResp_3_valid; // @[Cache.scala 175:22]
  wire  _T_24 = metaWay_0_tag == addr_tag; // @[Cache.scala 178:59]
  wire  _T_25 = metaWay_0_valid & _T_24; // @[Cache.scala 178:49]
  wire  _T_26 = _T_25 & io_in_valid; // @[Cache.scala 178:73]
  wire  _T_27 = metaWay_1_tag == addr_tag; // @[Cache.scala 178:59]
  wire  _T_28 = metaWay_1_valid & _T_27; // @[Cache.scala 178:49]
  wire  _T_29 = _T_28 & io_in_valid; // @[Cache.scala 178:73]
  wire  _T_30 = metaWay_2_tag == addr_tag; // @[Cache.scala 178:59]
  wire  _T_31 = metaWay_2_valid & _T_30; // @[Cache.scala 178:49]
  wire  _T_32 = _T_31 & io_in_valid; // @[Cache.scala 178:73]
  wire  _T_33 = metaWay_3_tag == addr_tag; // @[Cache.scala 178:59]
  wire  _T_34 = metaWay_3_valid & _T_33; // @[Cache.scala 178:49]
  wire  _T_35 = _T_34 & io_in_valid; // @[Cache.scala 178:73]
  wire [3:0] hitVec = {_T_35,_T_32,_T_29,_T_26}; // @[Cache.scala 178:90]
  reg [63:0] _T_39; // @[LFSR64.scala 25:23]
  wire  _T_42 = _T_39[0] ^ _T_39[1]; // @[LFSR64.scala 26:23]
  wire  _T_44 = _T_42 ^ _T_39[3]; // @[LFSR64.scala 26:33]
  wire  _T_46 = _T_44 ^ _T_39[4]; // @[LFSR64.scala 26:43]
  wire  _T_47 = _T_39 == 64'h0; // @[LFSR64.scala 28:24]
  wire [63:0] _T_49 = {_T_46,_T_39[63:1]}; // @[Cat.scala 29:58]
  wire [3:0] victimWaymask = 4'h1 << _T_39[1:0]; // @[Cache.scala 179:42]
  wire  _T_52 = ~metaWay_0_valid; // @[Cache.scala 181:45]
  wire  _T_53 = ~metaWay_1_valid; // @[Cache.scala 181:45]
  wire  _T_54 = ~metaWay_2_valid; // @[Cache.scala 181:45]
  wire  _T_55 = ~metaWay_3_valid; // @[Cache.scala 181:45]
  wire [3:0] invalidVec = {_T_55,_T_54,_T_53,_T_52}; // @[Cache.scala 181:56]
  wire  hasInvalidWay = |invalidVec; // @[Cache.scala 182:34]
  wire  _T_59 = invalidVec >= 4'h8; // @[Cache.scala 183:45]
  wire  _T_60 = invalidVec >= 4'h4; // @[Cache.scala 184:20]
  wire  _T_61 = invalidVec >= 4'h2; // @[Cache.scala 185:20]
  wire [1:0] _T_62 = _T_61 ? 2'h2 : 2'h1; // @[Cache.scala 185:8]
  wire [2:0] _T_63 = _T_60 ? 3'h4 : {{1'd0}, _T_62}; // @[Cache.scala 184:8]
  wire [3:0] refillInvalidWaymask = _T_59 ? 4'h8 : {{1'd0}, _T_63}; // @[Cache.scala 183:33]
  wire [3:0] _T_64 = hasInvalidWay ? refillInvalidWaymask : victimWaymask; // @[Cache.scala 188:49]
  wire [3:0] waymask = io_out_bits_hit ? hitVec : _T_64; // @[Cache.scala 188:20]
  wire [1:0] _T_69 = waymask[0] + waymask[1]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_71 = waymask[2] + waymask[3]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_73 = _T_69 + _T_71; // @[Bitwise.scala 47:55]
  wire  _T_75 = _T_73 > 3'h1; // @[Cache.scala 189:26]
  wire  _T_197 = io_in_valid & _T_75; // @[Cache.scala 196:24]
  wire  _T_198 = ~_T_197; // @[Cache.scala 196:10]
  wire  _T_200 = _T_198 | reset; // @[Cache.scala 196:9]
  wire  _T_201 = ~_T_200; // @[Cache.scala 196:9]
  wire  _T_202 = |hitVec; // @[Cache.scala 199:44]
  wire [31:0] _T_204 = io_in_bits_req_addr ^ 32'h30000000; // @[NutCore.scala 86:11]
  wire  _T_206 = _T_204[31:28] == 4'h0; // @[NutCore.scala 86:44]
  wire [31:0] _T_207 = io_in_bits_req_addr ^ 32'he0000000; // @[NutCore.scala 86:11]
  wire  _T_209 = _T_207[31:29] == 3'h0; // @[NutCore.scala 86:44]
  wire [9:0] _T_223 = {addr_index,addr_wordIndex}; // @[Cat.scala 29:58]
  wire  _T_224 = io_dataWriteBus_req_bits_setIdx == _T_223; // @[Cache.scala 205:30]
  wire  _T_225 = io_dataWriteBus_req_valid & _T_224; // @[Cache.scala 205:13]
  wire  isForwardData = io_in_valid & _T_225; // @[Cache.scala 204:35]
  reg  isForwardDataReg; // @[Cache.scala 207:33]
  wire  _GEN_8 = isForwardData | isForwardDataReg; // @[Cache.scala 208:24]
  reg [63:0] forwardDataReg_data_data; // @[Reg.scala 15:16]
  reg [3:0] forwardDataReg_waymask; // @[Reg.scala 15:16]
  wire  _T_232 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign io_in_ready = _T_14 | _T_232; // @[Cache.scala 216:15]
  assign io_out_valid = io_in_valid; // @[Cache.scala 215:16]
  assign io_out_bits_req_addr = io_in_bits_req_addr; // @[Cache.scala 214:19]
  assign io_out_bits_req_user = io_in_bits_req_user; // @[Cache.scala 214:19]
  assign io_out_bits_metas_0_tag = _T_16 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 198:21]
  assign io_out_bits_metas_0_valid = _T_16 | io_metaReadResp_0_valid; // @[Cache.scala 198:21]
  assign io_out_bits_metas_0_dirty = _T_16 ? _GEN_3 : io_metaReadResp_0_dirty; // @[Cache.scala 198:21]
  assign io_out_bits_metas_1_tag = _T_18 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 198:21]
  assign io_out_bits_metas_1_valid = _T_18 | io_metaReadResp_1_valid; // @[Cache.scala 198:21]
  assign io_out_bits_metas_1_dirty = _T_18 ? _GEN_3 : io_metaReadResp_1_dirty; // @[Cache.scala 198:21]
  assign io_out_bits_metas_2_tag = _T_20 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 198:21]
  assign io_out_bits_metas_2_valid = _T_20 | io_metaReadResp_2_valid; // @[Cache.scala 198:21]
  assign io_out_bits_metas_2_dirty = _T_20 ? _GEN_3 : io_metaReadResp_2_dirty; // @[Cache.scala 198:21]
  assign io_out_bits_metas_3_tag = _T_22 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 198:21]
  assign io_out_bits_metas_3_valid = _T_22 | io_metaReadResp_3_valid; // @[Cache.scala 198:21]
  assign io_out_bits_metas_3_dirty = _T_22 ? _GEN_3 : io_metaReadResp_3_dirty; // @[Cache.scala 198:21]
  assign io_out_bits_datas_0_data = io_dataReadResp_0_data; // @[Cache.scala 201:21]
  assign io_out_bits_datas_1_data = io_dataReadResp_1_data; // @[Cache.scala 201:21]
  assign io_out_bits_datas_2_data = io_dataReadResp_2_data; // @[Cache.scala 201:21]
  assign io_out_bits_datas_3_data = io_dataReadResp_3_data; // @[Cache.scala 201:21]
  assign io_out_bits_hit = io_in_valid & _T_202; // @[Cache.scala 199:19]
  assign io_out_bits_waymask = io_out_bits_hit ? hitVec : _T_64; // @[Cache.scala 200:23]
  assign io_out_bits_mmio = _T_206 | _T_209; // @[Cache.scala 202:20]
  assign io_out_bits_isForwardData = isForwardDataReg | isForwardData; // @[Cache.scala 211:29]
  assign io_out_bits_forwardData_data_data = isForwardData ? io_dataWriteBus_req_bits_data_data : forwardDataReg_data_data; // @[Cache.scala 212:27]
  assign io_out_bits_forwardData_waymask = isForwardData ? io_dataWriteBus_req_bits_waymask : forwardDataReg_waymask; // @[Cache.scala 212:27]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  isForwardMetaReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  forwardMetaReg_data_tag = _RAND_1[18:0];
  _RAND_2 = {1{`RANDOM}};
  forwardMetaReg_data_dirty = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  forwardMetaReg_waymask = _RAND_3[3:0];
  _RAND_4 = {2{`RANDOM}};
  _T_39 = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  isForwardDataReg = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  forwardDataReg_data_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  forwardDataReg_waymask = _RAND_7[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      isForwardMetaReg <= 1'h0;
    end else if (_T_15) begin
      isForwardMetaReg <= 1'h0;
    end else begin
      isForwardMetaReg <= _GEN_0;
    end
    if (isForwardMeta) begin
      forwardMetaReg_data_tag <= io_metaWriteBus_req_bits_data_tag;
    end
    if (isForwardMeta) begin
      forwardMetaReg_data_dirty <= io_metaWriteBus_req_bits_data_dirty;
    end
    if (isForwardMeta) begin
      forwardMetaReg_waymask <= io_metaWriteBus_req_bits_waymask;
    end
    if (reset) begin
      _T_39 <= 64'h1234567887654321;
    end else if (_T_47) begin
      _T_39 <= 64'h1;
    end else begin
      _T_39 <= _T_49;
    end
    if (reset) begin
      isForwardDataReg <= 1'h0;
    end else if (_T_15) begin
      isForwardDataReg <= 1'h0;
    end else begin
      isForwardDataReg <= _GEN_8;
    end
    if (isForwardData) begin
      forwardDataReg_data_data <= io_dataWriteBus_req_bits_data_data;
    end
    if (isForwardData) begin
      forwardDataReg_waymask <= io_dataWriteBus_req_bits_waymask;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_201) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Cache.scala:196 assert(!(io.in.valid && PopCount(waymask) > 1.U))\n"); // @[Cache.scala 196:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_201) begin
          $fatal; // @[Cache.scala 196:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Arbiter(
  input         io_in_0_valid,
  input  [6:0]  io_in_0_bits_setIdx,
  input  [18:0] io_in_0_bits_data_tag,
  input         io_in_0_bits_data_dirty,
  input  [3:0]  io_in_0_bits_waymask,
  input         io_in_1_valid,
  input  [6:0]  io_in_1_bits_setIdx,
  input  [18:0] io_in_1_bits_data_tag,
  input         io_in_1_bits_data_dirty,
  input  [3:0]  io_in_1_bits_waymask,
  output        io_out_valid,
  output [6:0]  io_out_bits_setIdx,
  output [18:0] io_out_bits_data_tag,
  output        io_out_bits_data_dirty,
  output [3:0]  io_out_bits_waymask
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  _T_2 = ~grant_1; // @[Arbiter.scala 135:19]
  assign io_out_valid = _T_2 | io_in_1_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_data_tag = io_in_0_valid ? io_in_0_bits_data_tag : io_in_1_bits_data_tag; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_data_dirty = io_in_0_valid ? io_in_0_bits_data_dirty : io_in_1_bits_data_dirty; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_waymask = io_in_0_valid ? io_in_0_bits_waymask : io_in_1_bits_waymask; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
endmodule
module Arbiter_1(
  input         io_in_0_valid,
  input  [9:0]  io_in_0_bits_setIdx,
  input  [63:0] io_in_0_bits_data_data,
  input  [3:0]  io_in_0_bits_waymask,
  input         io_in_1_valid,
  input  [9:0]  io_in_1_bits_setIdx,
  input  [63:0] io_in_1_bits_data_data,
  input  [3:0]  io_in_1_bits_waymask,
  output        io_out_valid,
  output [9:0]  io_out_bits_setIdx,
  output [63:0] io_out_bits_data_data,
  output [3:0]  io_out_bits_waymask
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  _T_2 = ~grant_1; // @[Arbiter.scala 135:19]
  assign io_out_valid = _T_2 | io_in_1_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_data_data = io_in_0_valid ? io_in_0_bits_data_data : io_in_1_bits_data_data; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_waymask = io_in_0_valid ? io_in_0_bits_waymask : io_in_1_bits_waymask; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
endmodule
module CacheStage3(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [86:0] io_in_bits_req_user,
  input  [18:0] io_in_bits_metas_0_tag,
  input         io_in_bits_metas_0_valid,
  input         io_in_bits_metas_0_dirty,
  input  [18:0] io_in_bits_metas_1_tag,
  input         io_in_bits_metas_1_valid,
  input         io_in_bits_metas_1_dirty,
  input  [18:0] io_in_bits_metas_2_tag,
  input         io_in_bits_metas_2_valid,
  input         io_in_bits_metas_2_dirty,
  input  [18:0] io_in_bits_metas_3_tag,
  input         io_in_bits_metas_3_valid,
  input         io_in_bits_metas_3_dirty,
  input  [63:0] io_in_bits_datas_0_data,
  input  [63:0] io_in_bits_datas_1_data,
  input  [63:0] io_in_bits_datas_2_data,
  input  [63:0] io_in_bits_datas_3_data,
  input         io_in_bits_hit,
  input  [3:0]  io_in_bits_waymask,
  input         io_in_bits_mmio,
  input         io_in_bits_isForwardData,
  input  [63:0] io_in_bits_forwardData_data_data,
  input  [3:0]  io_in_bits_forwardData_waymask,
  input         io_out_ready,
  output        io_out_valid,
  output [63:0] io_out_bits_rdata,
  output [86:0] io_out_bits_user,
  output        io_isFinish,
  input         io_flush,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [9:0]  io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data,
  output        io_dataWriteBus_req_valid,
  output [9:0]  io_dataWriteBus_req_bits_setIdx,
  output [63:0] io_dataWriteBus_req_bits_data_data,
  output [3:0]  io_dataWriteBus_req_bits_waymask,
  output        io_metaWriteBus_req_valid,
  output [6:0]  io_metaWriteBus_req_bits_setIdx,
  output [18:0] io_metaWriteBus_req_bits_data_tag,
  output        io_metaWriteBus_req_bits_data_dirty,
  output [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [31:0] io_mem_req_bits_addr,
  output [3:0]  io_mem_req_bits_cmd,
  output [63:0] io_mem_req_bits_wdata,
  output        io_mem_resp_ready,
  input         io_mem_resp_valid,
  input  [3:0]  io_mem_resp_bits_cmd,
  input  [63:0] io_mem_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  output        io_mmio_resp_ready,
  input         io_mmio_resp_valid,
  input  [63:0] io_mmio_resp_bits_rdata,
  output        io_cohResp_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
`endif // RANDOMIZE_REG_INIT
  wire  metaWriteArb_io_in_0_valid; // @[Cache.scala 241:28]
  wire [6:0] metaWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 241:28]
  wire [18:0] metaWriteArb_io_in_0_bits_data_tag; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_in_0_bits_data_dirty; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_in_0_bits_waymask; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_in_1_valid; // @[Cache.scala 241:28]
  wire [6:0] metaWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 241:28]
  wire [18:0] metaWriteArb_io_in_1_bits_data_tag; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_in_1_bits_data_dirty; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_in_1_bits_waymask; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_out_valid; // @[Cache.scala 241:28]
  wire [6:0] metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 241:28]
  wire [18:0] metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_out_bits_waymask; // @[Cache.scala 241:28]
  wire  dataWriteArb_io_in_0_valid; // @[Cache.scala 242:28]
  wire [9:0] dataWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 242:28]
  wire [63:0] dataWriteArb_io_in_0_bits_data_data; // @[Cache.scala 242:28]
  wire [3:0] dataWriteArb_io_in_0_bits_waymask; // @[Cache.scala 242:28]
  wire  dataWriteArb_io_in_1_valid; // @[Cache.scala 242:28]
  wire [9:0] dataWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 242:28]
  wire [63:0] dataWriteArb_io_in_1_bits_data_data; // @[Cache.scala 242:28]
  wire [3:0] dataWriteArb_io_in_1_bits_waymask; // @[Cache.scala 242:28]
  wire  dataWriteArb_io_out_valid; // @[Cache.scala 242:28]
  wire [9:0] dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 242:28]
  wire [63:0] dataWriteArb_io_out_bits_data_data; // @[Cache.scala 242:28]
  wire [3:0] dataWriteArb_io_out_bits_waymask; // @[Cache.scala 242:28]
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 245:31]
  wire [6:0] addr_index = io_in_bits_req_addr[12:6]; // @[Cache.scala 245:31]
  wire  mmio = io_in_valid & io_in_bits_mmio; // @[Cache.scala 246:26]
  wire  hit = io_in_valid & io_in_bits_hit; // @[Cache.scala 247:25]
  wire  _T_5 = ~io_in_bits_hit; // @[Cache.scala 248:29]
  wire  miss = io_in_valid & _T_5; // @[Cache.scala 248:26]
  wire [20:0] _T_14 = {io_in_bits_metas_0_tag,io_in_bits_metas_0_valid,io_in_bits_metas_0_dirty}; // @[Mux.scala 27:72]
  wire [20:0] _T_15 = io_in_bits_waymask[0] ? _T_14 : 21'h0; // @[Mux.scala 27:72]
  wire [20:0] _T_17 = {io_in_bits_metas_1_tag,io_in_bits_metas_1_valid,io_in_bits_metas_1_dirty}; // @[Mux.scala 27:72]
  wire [20:0] _T_18 = io_in_bits_waymask[1] ? _T_17 : 21'h0; // @[Mux.scala 27:72]
  wire [20:0] _T_20 = {io_in_bits_metas_2_tag,io_in_bits_metas_2_valid,io_in_bits_metas_2_dirty}; // @[Mux.scala 27:72]
  wire [20:0] _T_21 = io_in_bits_waymask[2] ? _T_20 : 21'h0; // @[Mux.scala 27:72]
  wire [20:0] _T_23 = {io_in_bits_metas_3_tag,io_in_bits_metas_3_valid,io_in_bits_metas_3_dirty}; // @[Mux.scala 27:72]
  wire [20:0] _T_24 = io_in_bits_waymask[3] ? _T_23 : 21'h0; // @[Mux.scala 27:72]
  wire [20:0] _T_25 = _T_15 | _T_18; // @[Mux.scala 27:72]
  wire [20:0] _T_26 = _T_25 | _T_21; // @[Mux.scala 27:72]
  wire [20:0] _T_27 = _T_26 | _T_24; // @[Mux.scala 27:72]
  wire [18:0] meta_tag = _T_27[20:2]; // @[Mux.scala 27:72]
  wire  _T_32 = mmio & hit; // @[Cache.scala 252:17]
  wire  _T_33 = ~_T_32; // @[Cache.scala 252:10]
  wire  _T_35 = _T_33 | reset; // @[Cache.scala 252:9]
  wire  _T_36 = ~_T_35; // @[Cache.scala 252:9]
  wire  _T_37 = io_in_bits_waymask == io_in_bits_forwardData_waymask; // @[Cache.scala 260:71]
  wire  useForwardData = io_in_bits_isForwardData & _T_37; // @[Cache.scala 260:49]
  wire [63:0] _T_42 = io_in_bits_waymask[0] ? io_in_bits_datas_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_43 = io_in_bits_waymask[1] ? io_in_bits_datas_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_44 = io_in_bits_waymask[2] ? io_in_bits_datas_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_45 = io_in_bits_waymask[3] ? io_in_bits_datas_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_46 = _T_42 | _T_43; // @[Mux.scala 27:72]
  wire [63:0] _T_47 = _T_46 | _T_44; // @[Mux.scala 27:72]
  wire [63:0] _T_48 = _T_47 | _T_45; // @[Mux.scala 27:72]
  wire [63:0] dataRead = useForwardData ? io_in_bits_forwardData_data_data : _T_48; // @[Cache.scala 262:21]
  wire  _T_86 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  reg [3:0] state; // @[Cache.scala 281:22]
  reg  needFlush; // @[Cache.scala 282:26]
  wire  _T_114 = state != 4'h0; // @[Cache.scala 284:28]
  wire  _T_115 = io_flush & _T_114; // @[Cache.scala 284:18]
  wire  _GEN_1 = _T_115 | needFlush; // @[Cache.scala 284:41]
  wire  _T_117 = _T_86 & needFlush; // @[Cache.scala 285:23]
  reg [2:0] value_1; // @[Counter.scala 29:33]
  reg [2:0] value_2; // @[Counter.scala 29:33]
  reg [1:0] state2; // @[Cache.scala 291:23]
  wire  _T_118 = state == 4'h3; // @[Cache.scala 293:39]
  wire  _T_119 = state == 4'h8; // @[Cache.scala 293:66]
  wire  _T_120 = _T_118 | _T_119; // @[Cache.scala 293:57]
  wire  _T_121 = state2 == 2'h0; // @[Cache.scala 293:92]
  wire [2:0] _T_124 = _T_119 ? value_1 : value_2; // @[Cache.scala 294:33]
  wire  _T_126 = state2 == 2'h1; // @[Cache.scala 295:60]
  reg [63:0] dataWay_0_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_1_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_2_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_3_data; // @[Reg.scala 15:16]
  wire [63:0] _T_131 = io_in_bits_waymask[0] ? dataWay_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_132 = io_in_bits_waymask[1] ? dataWay_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_133 = io_in_bits_waymask[2] ? dataWay_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_134 = io_in_bits_waymask[3] ? dataWay_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_135 = _T_131 | _T_132; // @[Mux.scala 27:72]
  wire [63:0] _T_136 = _T_135 | _T_133; // @[Mux.scala 27:72]
  wire  _T_141 = 2'h0 == state2; // @[Conditional.scala 37:30]
  wire  _T_142 = io_dataReadBus_req_ready & io_dataReadBus_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_143 = 2'h1 == state2; // @[Conditional.scala 37:30]
  wire  _T_144 = 2'h2 == state2; // @[Conditional.scala 37:30]
  wire  _T_145 = io_mem_req_ready & io_mem_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_147 = _T_145 | io_cohResp_valid; // @[Cache.scala 301:46]
  wire [31:0] raddr = {io_in_bits_req_addr[31:3],3'h0}; // @[Cat.scala 29:58]
  wire [31:0] waddr = {meta_tag,addr_index,6'h0}; // @[Cat.scala 29:58]
  wire  _T_152 = state == 4'h1; // @[Cache.scala 309:23]
  wire  _T_153 = value_2 == 3'h7; // @[Cache.scala 310:29]
  wire [2:0] _T_154 = _T_153 ? 3'h7 : 3'h3; // @[Cache.scala 310:8]
  wire [2:0] cmd = _T_152 ? 3'h2 : _T_154; // @[Cache.scala 309:16]
  wire  _T_160 = state2 == 2'h2; // @[Cache.scala 316:89]
  wire  _T_161 = _T_118 & _T_160; // @[Cache.scala 316:78]
  reg  afterFirstRead; // @[Cache.scala 323:31]
  reg  alreadyOutFire; // @[Reg.scala 27:20]
  wire  _GEN_12 = _T_86 | alreadyOutFire; // @[Reg.scala 28:19]
  wire  _T_165 = ~afterFirstRead; // @[Cache.scala 325:22]
  wire  _T_166 = io_mem_resp_ready & io_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_167 = _T_165 & _T_166; // @[Cache.scala 325:38]
  wire  _T_168 = state == 4'h2; // @[Cache.scala 325:70]
  wire  readingFirst = _T_167 & _T_168; // @[Cache.scala 325:60]
  wire  _T_170 = state == 4'h6; // @[Cache.scala 327:52]
  wire  _T_171 = mmio ? _T_170 : readingFirst; // @[Cache.scala 327:39]
  reg [63:0] inRdataRegDemand; // @[Reg.scala 15:16]
  wire  _T_172 = state == 4'h0; // @[Cache.scala 330:31]
  wire  _T_202 = 4'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_210 = miss | mmio; // @[Cache.scala 353:26]
  wire  _T_211 = ~io_flush; // @[Cache.scala 353:38]
  wire  _T_212 = _T_210 & _T_211; // @[Cache.scala 353:35]
  wire  _T_217 = 4'h5 == state; // @[Conditional.scala 37:30]
  wire  _T_218 = io_mmio_req_ready & io_mmio_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_219 = 4'h6 == state; // @[Conditional.scala 37:30]
  wire  _T_220 = io_mmio_resp_ready & io_mmio_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_221 = 4'h8 == state; // @[Conditional.scala 37:30]
  wire [2:0] _T_226 = value_1 + 3'h1; // @[Counter.scala 39:22]
  wire  _T_232 = 4'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_234 = 4'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_240 = io_mem_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire  _GEN_33 = _T_166 | afterFirstRead; // @[Cache.scala 372:33]
  wire  _T_241 = 4'h3 == state; // @[Conditional.scala 37:30]
  wire [2:0] _T_245 = value_2 + 3'h1; // @[Counter.scala 39:22]
  wire  _T_246 = io_mem_req_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_248 = _T_246 & _T_145; // @[Cache.scala 382:43]
  wire  _T_249 = 4'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_251 = 4'h7 == state; // @[Conditional.scala 37:30]
  wire  _T_253 = _T_86 | needFlush; // @[Cache.scala 386:44]
  wire  _T_254 = _T_253 | alreadyOutFire; // @[Cache.scala 386:57]
  wire  dataRefillWriteBus_req_valid = _T_168 & _T_166; // @[Cache.scala 391:39]
  wire  _T_293 = state == 4'h7; // @[Cache.scala 433:48]
  wire  _T_310 = ~alreadyOutFire; // @[Cache.scala 434:110]
  wire  _T_311 = afterFirstRead & _T_310; // @[Cache.scala 434:107]
  wire  _T_312 = mmio ? _T_293 : _T_311; // @[Cache.scala 434:45]
  wire  _T_313 = hit | _T_312; // @[Cache.scala 434:28]
  wire  _T_329 = _T_293 & _GEN_12; // @[Cache.scala 442:70]
  wire  _T_335 = io_out_ready & _T_172; // @[Cache.scala 445:31]
  wire  _T_336 = ~miss; // @[Cache.scala 445:73]
  Arbiter metaWriteArb ( // @[Cache.scala 241:28]
    .io_in_0_valid(metaWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(metaWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_tag(metaWriteArb_io_in_0_bits_data_tag),
    .io_in_0_bits_data_dirty(metaWriteArb_io_in_0_bits_data_dirty),
    .io_in_0_bits_waymask(metaWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(metaWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(metaWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_tag(metaWriteArb_io_in_1_bits_data_tag),
    .io_in_1_bits_data_dirty(metaWriteArb_io_in_1_bits_data_dirty),
    .io_in_1_bits_waymask(metaWriteArb_io_in_1_bits_waymask),
    .io_out_valid(metaWriteArb_io_out_valid),
    .io_out_bits_setIdx(metaWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_tag(metaWriteArb_io_out_bits_data_tag),
    .io_out_bits_data_dirty(metaWriteArb_io_out_bits_data_dirty),
    .io_out_bits_waymask(metaWriteArb_io_out_bits_waymask)
  );
  Arbiter_1 dataWriteArb ( // @[Cache.scala 242:28]
    .io_in_0_valid(dataWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(dataWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_data(dataWriteArb_io_in_0_bits_data_data),
    .io_in_0_bits_waymask(dataWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(dataWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(dataWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_data(dataWriteArb_io_in_1_bits_data_data),
    .io_in_1_bits_waymask(dataWriteArb_io_in_1_bits_waymask),
    .io_out_valid(dataWriteArb_io_out_valid),
    .io_out_bits_setIdx(dataWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_data(dataWriteArb_io_out_bits_data_data),
    .io_out_bits_waymask(dataWriteArb_io_out_bits_waymask)
  );
  assign io_in_ready = _T_335 & _T_336; // @[Cache.scala 445:15]
  assign io_out_valid = io_in_valid & _T_313; // @[Cache.scala 432:16]
  assign io_out_bits_rdata = hit ? dataRead : inRdataRegDemand; // @[Cache.scala 426:23]
  assign io_out_bits_user = io_in_bits_req_user; // @[Cache.scala 429:56]
  assign io_isFinish = hit ? _T_86 : _T_329; // @[Cache.scala 441:15]
  assign io_dataReadBus_req_valid = _T_120 & _T_121; // @[SRAMTemplate.scala 53:20]
  assign io_dataReadBus_req_bits_setIdx = {addr_index,_T_124}; // @[SRAMTemplate.scala 26:17]
  assign io_dataWriteBus_req_valid = dataWriteArb_io_out_valid; // @[Cache.scala 396:23]
  assign io_dataWriteBus_req_bits_setIdx = dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 396:23]
  assign io_dataWriteBus_req_bits_data_data = dataWriteArb_io_out_bits_data_data; // @[Cache.scala 396:23]
  assign io_dataWriteBus_req_bits_waymask = dataWriteArb_io_out_bits_waymask; // @[Cache.scala 396:23]
  assign io_metaWriteBus_req_valid = metaWriteArb_io_out_valid; // @[Cache.scala 406:23]
  assign io_metaWriteBus_req_bits_setIdx = metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 406:23]
  assign io_metaWriteBus_req_bits_data_tag = metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 406:23]
  assign io_metaWriteBus_req_bits_data_dirty = metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 406:23]
  assign io_metaWriteBus_req_bits_waymask = metaWriteArb_io_out_bits_waymask; // @[Cache.scala 406:23]
  assign io_mem_req_valid = _T_152 | _T_161; // @[Cache.scala 316:20]
  assign io_mem_req_bits_addr = _T_152 ? raddr : waddr; // @[SimpleBus.scala 64:15]
  assign io_mem_req_bits_cmd = {{1'd0}, cmd}; // @[SimpleBus.scala 65:14]
  assign io_mem_req_bits_wdata = _T_136 | _T_134; // @[SimpleBus.scala 67:16]
  assign io_mem_resp_ready = 1'h1; // @[Cache.scala 315:21]
  assign io_mmio_req_valid = state == 4'h5; // @[Cache.scala 321:21]
  assign io_mmio_req_bits_addr = io_in_bits_req_addr; // @[Cache.scala 319:20]
  assign io_mmio_resp_ready = 1'h1; // @[Cache.scala 320:22]
  assign io_cohResp_valid = _T_119 & _T_160; // @[Cache.scala 330:20]
  assign metaWriteArb_io_in_0_valid = 1'h0; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_0_bits_setIdx = io_in_bits_req_addr[12:6]; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_0_bits_data_tag = _T_27[20:2]; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_0_bits_data_dirty = 1'h0; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_1_valid = dataRefillWriteBus_req_valid & _T_240; // @[Cache.scala 405:25]
  assign metaWriteArb_io_in_1_bits_setIdx = io_in_bits_req_addr[12:6]; // @[Cache.scala 405:25]
  assign metaWriteArb_io_in_1_bits_data_tag = io_in_bits_req_addr[31:13]; // @[Cache.scala 405:25]
  assign metaWriteArb_io_in_1_bits_data_dirty = 1'h0; // @[Cache.scala 405:25]
  assign metaWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 405:25]
  assign dataWriteArb_io_in_0_valid = 1'h0; // @[Cache.scala 394:25]
  assign dataWriteArb_io_in_0_bits_setIdx = {addr_index,addr_wordIndex}; // @[Cache.scala 394:25]
  assign dataWriteArb_io_in_0_bits_data_data = useForwardData ? io_in_bits_forwardData_data_data : _T_48; // @[Cache.scala 394:25]
  assign dataWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 394:25]
  assign dataWriteArb_io_in_1_valid = _T_168 & _T_166; // @[Cache.scala 395:25]
  assign dataWriteArb_io_in_1_bits_setIdx = {addr_index,value_1}; // @[Cache.scala 395:25]
  assign dataWriteArb_io_in_1_bits_data_data = io_mem_resp_bits_rdata; // @[Cache.scala 395:25]
  assign dataWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 395:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[3:0];
  _RAND_1 = {1{`RANDOM}};
  needFlush = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  value_2 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  state2 = _RAND_4[1:0];
  _RAND_5 = {2{`RANDOM}};
  dataWay_0_data = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  dataWay_1_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  dataWay_2_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  dataWay_3_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  afterFirstRead = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  alreadyOutFire = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  inRdataRegDemand = _RAND_11[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 4'h0;
    end else if (_T_202) begin
      if (_T_212) begin
        if (mmio) begin
          state <= 4'h5;
        end else begin
          state <= 4'h1;
        end
      end
    end else if (_T_217) begin
      if (_T_218) begin
        state <= 4'h6;
      end
    end else if (_T_219) begin
      if (_T_220) begin
        state <= 4'h7;
      end
    end else if (!(_T_221)) begin
      if (_T_232) begin
        if (_T_145) begin
          state <= 4'h2;
        end
      end else if (_T_234) begin
        if (_T_166) begin
          if (_T_240) begin
            state <= 4'h7;
          end
        end
      end else if (_T_241) begin
        if (_T_248) begin
          state <= 4'h4;
        end
      end else if (_T_249) begin
        if (_T_166) begin
          state <= 4'h1;
        end
      end else if (_T_251) begin
        if (_T_254) begin
          state <= 4'h0;
        end
      end
    end
    if (reset) begin
      needFlush <= 1'h0;
    end else if (_T_117) begin
      needFlush <= 1'h0;
    end else begin
      needFlush <= _GEN_1;
    end
    if (reset) begin
      value_1 <= 3'h0;
    end else if (!(_T_202)) begin
      if (!(_T_217)) begin
        if (!(_T_219)) begin
          if (_T_221) begin
            if (io_cohResp_valid) begin
              value_1 <= _T_226;
            end
          end else if (_T_232) begin
            if (_T_145) begin
              value_1 <= addr_wordIndex;
            end
          end else if (_T_234) begin
            if (_T_166) begin
              value_1 <= _T_226;
            end
          end
        end
      end
    end
    if (reset) begin
      value_2 <= 3'h0;
    end else if (!(_T_202)) begin
      if (!(_T_217)) begin
        if (!(_T_219)) begin
          if (!(_T_221)) begin
            if (!(_T_232)) begin
              if (!(_T_234)) begin
                if (_T_241) begin
                  if (_T_145) begin
                    value_2 <= _T_245;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      state2 <= 2'h0;
    end else if (_T_141) begin
      if (_T_142) begin
        state2 <= 2'h1;
      end
    end else if (_T_143) begin
      state2 <= 2'h2;
    end else if (_T_144) begin
      if (_T_147) begin
        state2 <= 2'h0;
      end
    end
    if (_T_126) begin
      dataWay_0_data <= io_dataReadBus_resp_data_0_data;
    end
    if (_T_126) begin
      dataWay_1_data <= io_dataReadBus_resp_data_1_data;
    end
    if (_T_126) begin
      dataWay_2_data <= io_dataReadBus_resp_data_2_data;
    end
    if (_T_126) begin
      dataWay_3_data <= io_dataReadBus_resp_data_3_data;
    end
    if (reset) begin
      afterFirstRead <= 1'h0;
    end else if (_T_202) begin
      afterFirstRead <= 1'h0;
    end else if (!(_T_217)) begin
      if (!(_T_219)) begin
        if (!(_T_221)) begin
          if (!(_T_232)) begin
            if (_T_234) begin
              afterFirstRead <= _GEN_33;
            end
          end
        end
      end
    end
    if (reset) begin
      alreadyOutFire <= 1'h0;
    end else if (_T_202) begin
      alreadyOutFire <= 1'h0;
    end else begin
      alreadyOutFire <= _GEN_12;
    end
    if (_T_171) begin
      if (mmio) begin
        inRdataRegDemand <= io_mmio_resp_bits_rdata;
      end else begin
        inRdataRegDemand <= io_mem_resp_bits_rdata;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_36) begin
          $fwrite(32'h80000002,"Assertion failed: MMIO request should not hit in cache\n    at Cache.scala:252 assert(!(mmio && hit), \"MMIO request should not hit in cache\")\n"); // @[Cache.scala 252:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_36) begin
          $fatal; // @[Cache.scala 252:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module SRAMTemplate_1(
  input         clock,
  input         reset,
  output        io_rreq_ready,
  input         io_rreq_valid,
  input  [6:0]  io_rreq_bits_setIdx,
  output [18:0] io_rresp_data_0_tag,
  output        io_rresp_data_0_valid,
  output        io_rresp_data_0_dirty,
  output [18:0] io_rresp_data_1_tag,
  output        io_rresp_data_1_valid,
  output        io_rresp_data_1_dirty,
  output [18:0] io_rresp_data_2_tag,
  output        io_rresp_data_2_valid,
  output        io_rresp_data_2_dirty,
  output [18:0] io_rresp_data_3_tag,
  output        io_rresp_data_3_valid,
  output        io_rresp_data_3_dirty,
  input         io_wreq_valid,
  input  [6:0]  io_wreq_bits_setIdx,
  input  [18:0] io_wreq_bits_data_tag,
  input         io_wreq_bits_data_dirty,
  input  [3:0]  io_wreq_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire [6:0] array_RW0_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_en; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_clk; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmode; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_RW0_wdata_0; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_RW0_wdata_1; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_RW0_wdata_2; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_RW0_wdata_3; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_RW0_rdata_0; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_RW0_rdata_1; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_RW0_rdata_2; // @[SRAMTemplate.scala 76:26]
  wire [20:0] array_RW0_rdata_3; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_0; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_1; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_2; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_3; // @[SRAMTemplate.scala 76:26]
  reg  resetState; // @[SRAMTemplate.scala 80:30]
  reg [6:0] resetSet; // @[Counter.scala 29:33]
  wire  _T_3 = resetSet == 7'h7f; // @[Counter.scala 38:24]
  wire [6:0] _T_5 = resetSet + 7'h1; // @[Counter.scala 39:22]
  wire  _GEN_1 = resetState & _T_3; // @[Counter.scala 67:17]
  wire  _GEN_2 = _GEN_1 ? 1'h0 : resetState; // @[SRAMTemplate.scala 82:24]
  wire  wen = io_wreq_valid | resetState; // @[SRAMTemplate.scala 88:52]
  wire  _T_6 = ~wen; // @[SRAMTemplate.scala 89:41]
  wire  realRen = io_rreq_valid & _T_6; // @[SRAMTemplate.scala 89:38]
  wire [6:0] setIdx = resetState ? resetSet : io_wreq_bits_setIdx; // @[SRAMTemplate.scala 91:19]
  wire [20:0] _T_9 = {io_wreq_bits_data_tag,1'h1,io_wreq_bits_data_dirty}; // @[SRAMTemplate.scala 92:78]
  wire [3:0] waymask = resetState ? 4'hf : io_wreq_bits_waymask; // @[SRAMTemplate.scala 93:20]
  wire [20:0] _T_22 = array_RW0_rdata_0;
  wire [20:0] _T_26 = array_RW0_rdata_1;
  wire [20:0] _T_30 = array_RW0_rdata_2;
  wire [20:0] _T_34 = array_RW0_rdata_3;
  wire  _T_39 = ~resetState; // @[SRAMTemplate.scala 101:21]
  array_0 array ( // @[SRAMTemplate.scala 76:26]
    .RW0_addr(array_RW0_addr),
    .RW0_en(array_RW0_en),
    .RW0_clk(array_RW0_clk),
    .RW0_wmode(array_RW0_wmode),
    .RW0_wdata_0(array_RW0_wdata_0),
    .RW0_wdata_1(array_RW0_wdata_1),
    .RW0_wdata_2(array_RW0_wdata_2),
    .RW0_wdata_3(array_RW0_wdata_3),
    .RW0_rdata_0(array_RW0_rdata_0),
    .RW0_rdata_1(array_RW0_rdata_1),
    .RW0_rdata_2(array_RW0_rdata_2),
    .RW0_rdata_3(array_RW0_rdata_3),
    .RW0_wmask_0(array_RW0_wmask_0),
    .RW0_wmask_1(array_RW0_wmask_1),
    .RW0_wmask_2(array_RW0_wmask_2),
    .RW0_wmask_3(array_RW0_wmask_3)
  );
  assign io_rreq_ready = _T_39 & _T_6; // @[SRAMTemplate.scala 101:18]
  assign io_rresp_data_0_tag = _T_22[20:2]; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_0_valid = _T_22[1]; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_0_dirty = _T_22[0]; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_1_tag = _T_26[20:2]; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_1_valid = _T_26[1]; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_1_dirty = _T_26[0]; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_2_tag = _T_30[20:2]; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_2_valid = _T_30[1]; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_2_dirty = _T_30[0]; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_3_tag = _T_34[20:2]; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_3_valid = _T_34[1]; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_3_dirty = _T_34[0]; // @[SRAMTemplate.scala 99:18]
  assign array_RW0_wdata_0 = resetState ? 21'h0 : _T_9;
  assign array_RW0_wdata_1 = resetState ? 21'h0 : _T_9;
  assign array_RW0_wdata_2 = resetState ? 21'h0 : _T_9;
  assign array_RW0_wdata_3 = resetState ? 21'h0 : _T_9;
  assign array_RW0_wmask_0 = waymask[0];
  assign array_RW0_wmask_1 = waymask[1];
  assign array_RW0_wmask_2 = waymask[2];
  assign array_RW0_wmask_3 = waymask[3];
  assign array_RW0_wmode = io_wreq_valid | resetState;
  assign array_RW0_clk = clock;
  assign array_RW0_en = realRen | wen;
  assign array_RW0_addr = wen ? setIdx : io_rreq_bits_setIdx;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  resetState = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  resetSet = _RAND_1[6:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    resetState <= reset | _GEN_2;
    if (reset) begin
      resetSet <= 7'h0;
    end else if (resetState) begin
      resetSet <= _T_5;
    end
  end
endmodule
module Arbiter_2(
  output       io_in_0_ready,
  input        io_in_0_valid,
  input  [6:0] io_in_0_bits_setIdx,
  input        io_out_ready,
  output       io_out_valid,
  output [6:0] io_out_bits_setIdx
);
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = io_in_0_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_setIdx = io_in_0_bits_setIdx; // @[Arbiter.scala 124:15]
endmodule
module SRAMTemplateWithArbiter(
  input         clock,
  input         reset,
  output        io_r0_req_ready,
  input         io_r0_req_valid,
  input  [6:0]  io_r0_req_bits_setIdx,
  output [18:0] io_r0_resp_data_0_tag,
  output        io_r0_resp_data_0_valid,
  output        io_r0_resp_data_0_dirty,
  output [18:0] io_r0_resp_data_1_tag,
  output        io_r0_resp_data_1_valid,
  output        io_r0_resp_data_1_dirty,
  output [18:0] io_r0_resp_data_2_tag,
  output        io_r0_resp_data_2_valid,
  output        io_r0_resp_data_2_dirty,
  output [18:0] io_r0_resp_data_3_tag,
  output        io_r0_resp_data_3_valid,
  output        io_r0_resp_data_3_dirty,
  input         io_wreq_valid,
  input  [6:0]  io_wreq_bits_setIdx,
  input  [18:0] io_wreq_bits_data_tag,
  input         io_wreq_bits_data_dirty,
  input  [3:0]  io_wreq_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  ram_clock; // @[SRAMTemplate.scala 121:19]
  wire  ram_reset; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rreq_ready; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rreq_valid; // @[SRAMTemplate.scala 121:19]
  wire [6:0] ram_io_rreq_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [18:0] ram_io_rresp_data_0_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_0_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_0_dirty; // @[SRAMTemplate.scala 121:19]
  wire [18:0] ram_io_rresp_data_1_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_1_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_1_dirty; // @[SRAMTemplate.scala 121:19]
  wire [18:0] ram_io_rresp_data_2_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_2_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_2_dirty; // @[SRAMTemplate.scala 121:19]
  wire [18:0] ram_io_rresp_data_3_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_3_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_3_dirty; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_wreq_valid; // @[SRAMTemplate.scala 121:19]
  wire [6:0] ram_io_wreq_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [18:0] ram_io_wreq_bits_data_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_wreq_bits_data_dirty; // @[SRAMTemplate.scala 121:19]
  wire [3:0] ram_io_wreq_bits_waymask; // @[SRAMTemplate.scala 121:19]
  wire  readArb_io_in_0_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_0_valid; // @[SRAMTemplate.scala 124:23]
  wire [6:0] readArb_io_in_0_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_valid; // @[SRAMTemplate.scala 124:23]
  wire [6:0] readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  reg  _T_1; // @[SRAMTemplate.scala 130:58]
  reg [18:0] _T_3_0_tag; // @[Reg.scala 27:20]
  reg  _T_3_0_valid; // @[Reg.scala 27:20]
  reg  _T_3_0_dirty; // @[Reg.scala 27:20]
  reg [18:0] _T_3_1_tag; // @[Reg.scala 27:20]
  reg  _T_3_1_valid; // @[Reg.scala 27:20]
  reg  _T_3_1_dirty; // @[Reg.scala 27:20]
  reg [18:0] _T_3_2_tag; // @[Reg.scala 27:20]
  reg  _T_3_2_valid; // @[Reg.scala 27:20]
  reg  _T_3_2_dirty; // @[Reg.scala 27:20]
  reg [18:0] _T_3_3_tag; // @[Reg.scala 27:20]
  reg  _T_3_3_valid; // @[Reg.scala 27:20]
  reg  _T_3_3_dirty; // @[Reg.scala 27:20]
  SRAMTemplate_1 ram ( // @[SRAMTemplate.scala 121:19]
    .clock(ram_clock),
    .reset(ram_reset),
    .io_rreq_ready(ram_io_rreq_ready),
    .io_rreq_valid(ram_io_rreq_valid),
    .io_rreq_bits_setIdx(ram_io_rreq_bits_setIdx),
    .io_rresp_data_0_tag(ram_io_rresp_data_0_tag),
    .io_rresp_data_0_valid(ram_io_rresp_data_0_valid),
    .io_rresp_data_0_dirty(ram_io_rresp_data_0_dirty),
    .io_rresp_data_1_tag(ram_io_rresp_data_1_tag),
    .io_rresp_data_1_valid(ram_io_rresp_data_1_valid),
    .io_rresp_data_1_dirty(ram_io_rresp_data_1_dirty),
    .io_rresp_data_2_tag(ram_io_rresp_data_2_tag),
    .io_rresp_data_2_valid(ram_io_rresp_data_2_valid),
    .io_rresp_data_2_dirty(ram_io_rresp_data_2_dirty),
    .io_rresp_data_3_tag(ram_io_rresp_data_3_tag),
    .io_rresp_data_3_valid(ram_io_rresp_data_3_valid),
    .io_rresp_data_3_dirty(ram_io_rresp_data_3_dirty),
    .io_wreq_valid(ram_io_wreq_valid),
    .io_wreq_bits_setIdx(ram_io_wreq_bits_setIdx),
    .io_wreq_bits_data_tag(ram_io_wreq_bits_data_tag),
    .io_wreq_bits_data_dirty(ram_io_wreq_bits_data_dirty),
    .io_wreq_bits_waymask(ram_io_wreq_bits_waymask)
  );
  Arbiter_2 readArb ( // @[SRAMTemplate.scala 124:23]
    .io_in_0_ready(readArb_io_in_0_ready),
    .io_in_0_valid(readArb_io_in_0_valid),
    .io_in_0_bits_setIdx(readArb_io_in_0_bits_setIdx),
    .io_out_ready(readArb_io_out_ready),
    .io_out_valid(readArb_io_out_valid),
    .io_out_bits_setIdx(readArb_io_out_bits_setIdx)
  );
  assign io_r0_req_ready = readArb_io_in_0_ready; // @[SRAMTemplate.scala 125:17]
  assign io_r0_resp_data_0_tag = _T_1 ? ram_io_rresp_data_0_tag : _T_3_0_tag; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_0_valid = _T_1 ? ram_io_rresp_data_0_valid : _T_3_0_valid; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_0_dirty = _T_1 ? ram_io_rresp_data_0_dirty : _T_3_0_dirty; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_1_tag = _T_1 ? ram_io_rresp_data_1_tag : _T_3_1_tag; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_1_valid = _T_1 ? ram_io_rresp_data_1_valid : _T_3_1_valid; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_1_dirty = _T_1 ? ram_io_rresp_data_1_dirty : _T_3_1_dirty; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_2_tag = _T_1 ? ram_io_rresp_data_2_tag : _T_3_2_tag; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_2_valid = _T_1 ? ram_io_rresp_data_2_valid : _T_3_2_valid; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_2_dirty = _T_1 ? ram_io_rresp_data_2_dirty : _T_3_2_dirty; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_3_tag = _T_1 ? ram_io_rresp_data_3_tag : _T_3_3_tag; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_3_valid = _T_1 ? ram_io_rresp_data_3_valid : _T_3_3_valid; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_3_dirty = _T_1 ? ram_io_rresp_data_3_dirty : _T_3_3_dirty; // @[SRAMTemplate.scala 130:17]
  assign ram_clock = clock;
  assign ram_reset = reset;
  assign ram_io_rreq_valid = readArb_io_out_valid; // @[SRAMTemplate.scala 126:16]
  assign ram_io_rreq_bits_setIdx = readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 126:16]
  assign ram_io_wreq_valid = io_wreq_valid; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_setIdx = io_wreq_bits_setIdx; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_data_tag = io_wreq_bits_data_tag; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_data_dirty = io_wreq_bits_data_dirty; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_waymask = io_wreq_bits_waymask; // @[SRAMTemplate.scala 122:12]
  assign readArb_io_in_0_valid = io_r0_req_valid; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_0_bits_setIdx = io_r0_req_bits_setIdx; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_out_ready = ram_io_rreq_ready; // @[SRAMTemplate.scala 126:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _T_3_0_tag = _RAND_1[18:0];
  _RAND_2 = {1{`RANDOM}};
  _T_3_0_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _T_3_0_dirty = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_3_1_tag = _RAND_4[18:0];
  _RAND_5 = {1{`RANDOM}};
  _T_3_1_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_3_1_dirty = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_3_2_tag = _RAND_7[18:0];
  _RAND_8 = {1{`RANDOM}};
  _T_3_2_valid = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _T_3_2_dirty = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _T_3_3_tag = _RAND_10[18:0];
  _RAND_11 = {1{`RANDOM}};
  _T_3_3_valid = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _T_3_3_dirty = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_1 <= io_r0_req_ready & io_r0_req_valid;
    if (reset) begin
      _T_3_0_tag <= 19'h0;
    end else if (_T_1) begin
      _T_3_0_tag <= ram_io_rresp_data_0_tag;
    end
    if (reset) begin
      _T_3_0_valid <= 1'h0;
    end else if (_T_1) begin
      _T_3_0_valid <= ram_io_rresp_data_0_valid;
    end
    if (reset) begin
      _T_3_0_dirty <= 1'h0;
    end else if (_T_1) begin
      _T_3_0_dirty <= ram_io_rresp_data_0_dirty;
    end
    if (reset) begin
      _T_3_1_tag <= 19'h0;
    end else if (_T_1) begin
      _T_3_1_tag <= ram_io_rresp_data_1_tag;
    end
    if (reset) begin
      _T_3_1_valid <= 1'h0;
    end else if (_T_1) begin
      _T_3_1_valid <= ram_io_rresp_data_1_valid;
    end
    if (reset) begin
      _T_3_1_dirty <= 1'h0;
    end else if (_T_1) begin
      _T_3_1_dirty <= ram_io_rresp_data_1_dirty;
    end
    if (reset) begin
      _T_3_2_tag <= 19'h0;
    end else if (_T_1) begin
      _T_3_2_tag <= ram_io_rresp_data_2_tag;
    end
    if (reset) begin
      _T_3_2_valid <= 1'h0;
    end else if (_T_1) begin
      _T_3_2_valid <= ram_io_rresp_data_2_valid;
    end
    if (reset) begin
      _T_3_2_dirty <= 1'h0;
    end else if (_T_1) begin
      _T_3_2_dirty <= ram_io_rresp_data_2_dirty;
    end
    if (reset) begin
      _T_3_3_tag <= 19'h0;
    end else if (_T_1) begin
      _T_3_3_tag <= ram_io_rresp_data_3_tag;
    end
    if (reset) begin
      _T_3_3_valid <= 1'h0;
    end else if (_T_1) begin
      _T_3_3_valid <= ram_io_rresp_data_3_valid;
    end
    if (reset) begin
      _T_3_3_dirty <= 1'h0;
    end else if (_T_1) begin
      _T_3_3_dirty <= ram_io_rresp_data_3_dirty;
    end
  end
endmodule
module SRAMTemplate_2(
  input         clock,
  output        io_rreq_ready,
  input         io_rreq_valid,
  input  [9:0]  io_rreq_bits_setIdx,
  output [63:0] io_rresp_data_0_data,
  output [63:0] io_rresp_data_1_data,
  output [63:0] io_rresp_data_2_data,
  output [63:0] io_rresp_data_3_data,
  input         io_wreq_valid,
  input  [9:0]  io_wreq_bits_setIdx,
  input  [63:0] io_wreq_bits_data_data,
  input  [3:0]  io_wreq_bits_waymask
);
  wire [9:0] array_RW0_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_en; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_clk; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmode; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_wdata_0; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_wdata_1; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_wdata_2; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_wdata_3; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_rdata_0; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_rdata_1; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_rdata_2; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_rdata_3; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_0; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_1; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_2; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_3; // @[SRAMTemplate.scala 76:26]
  wire  _T = ~io_wreq_valid; // @[SRAMTemplate.scala 89:41]
  wire  realRen = io_rreq_valid & _T; // @[SRAMTemplate.scala 89:38]
  array_1 array ( // @[SRAMTemplate.scala 76:26]
    .RW0_addr(array_RW0_addr),
    .RW0_en(array_RW0_en),
    .RW0_clk(array_RW0_clk),
    .RW0_wmode(array_RW0_wmode),
    .RW0_wdata_0(array_RW0_wdata_0),
    .RW0_wdata_1(array_RW0_wdata_1),
    .RW0_wdata_2(array_RW0_wdata_2),
    .RW0_wdata_3(array_RW0_wdata_3),
    .RW0_rdata_0(array_RW0_rdata_0),
    .RW0_rdata_1(array_RW0_rdata_1),
    .RW0_rdata_2(array_RW0_rdata_2),
    .RW0_rdata_3(array_RW0_rdata_3),
    .RW0_wmask_0(array_RW0_wmask_0),
    .RW0_wmask_1(array_RW0_wmask_1),
    .RW0_wmask_2(array_RW0_wmask_2),
    .RW0_wmask_3(array_RW0_wmask_3)
  );
  assign io_rreq_ready = ~io_wreq_valid; // @[SRAMTemplate.scala 101:18]
  assign io_rresp_data_0_data = array_RW0_rdata_0; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_1_data = array_RW0_rdata_1; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_2_data = array_RW0_rdata_2; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_3_data = array_RW0_rdata_3; // @[SRAMTemplate.scala 99:18]
  assign array_RW0_wdata_0 = io_wreq_bits_data_data;
  assign array_RW0_wdata_1 = io_wreq_bits_data_data;
  assign array_RW0_wdata_2 = io_wreq_bits_data_data;
  assign array_RW0_wdata_3 = io_wreq_bits_data_data;
  assign array_RW0_wmask_0 = io_wreq_bits_waymask[0];
  assign array_RW0_wmask_1 = io_wreq_bits_waymask[1];
  assign array_RW0_wmask_2 = io_wreq_bits_waymask[2];
  assign array_RW0_wmask_3 = io_wreq_bits_waymask[3];
  assign array_RW0_wmode = io_wreq_valid;
  assign array_RW0_clk = clock;
  assign array_RW0_en = realRen | io_wreq_valid;
  assign array_RW0_addr = io_wreq_valid ? io_wreq_bits_setIdx : io_rreq_bits_setIdx;
endmodule
module Arbiter_3(
  output       io_in_0_ready,
  input        io_in_0_valid,
  input  [9:0] io_in_0_bits_setIdx,
  output       io_in_1_ready,
  input        io_in_1_valid,
  input  [9:0] io_in_1_bits_setIdx,
  input        io_out_ready,
  output       io_out_valid,
  output [9:0] io_out_bits_setIdx
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  _T_2 = ~grant_1; // @[Arbiter.scala 135:19]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = _T_2 | io_in_1_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
endmodule
module SRAMTemplateWithArbiter_1(
  input         clock,
  input         reset,
  output        io_r0_req_ready,
  input         io_r0_req_valid,
  input  [9:0]  io_r0_req_bits_setIdx,
  output [63:0] io_r0_resp_data_0_data,
  output [63:0] io_r0_resp_data_1_data,
  output [63:0] io_r0_resp_data_2_data,
  output [63:0] io_r0_resp_data_3_data,
  output        io_r1_req_ready,
  input         io_r1_req_valid,
  input  [9:0]  io_r1_req_bits_setIdx,
  output [63:0] io_r1_resp_data_0_data,
  output [63:0] io_r1_resp_data_1_data,
  output [63:0] io_r1_resp_data_2_data,
  output [63:0] io_r1_resp_data_3_data,
  input         io_wreq_valid,
  input  [9:0]  io_wreq_bits_setIdx,
  input  [63:0] io_wreq_bits_data_data,
  input  [3:0]  io_wreq_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  ram_clock; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rreq_ready; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rreq_valid; // @[SRAMTemplate.scala 121:19]
  wire [9:0] ram_io_rreq_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_rresp_data_0_data; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_rresp_data_1_data; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_rresp_data_2_data; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_rresp_data_3_data; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_wreq_valid; // @[SRAMTemplate.scala 121:19]
  wire [9:0] ram_io_wreq_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_wreq_bits_data_data; // @[SRAMTemplate.scala 121:19]
  wire [3:0] ram_io_wreq_bits_waymask; // @[SRAMTemplate.scala 121:19]
  wire  readArb_io_in_0_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_0_valid; // @[SRAMTemplate.scala 124:23]
  wire [9:0] readArb_io_in_0_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_1_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_1_valid; // @[SRAMTemplate.scala 124:23]
  wire [9:0] readArb_io_in_1_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_valid; // @[SRAMTemplate.scala 124:23]
  wire [9:0] readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  reg  _T_1; // @[SRAMTemplate.scala 130:58]
  reg [63:0] _T_3_0_data; // @[Reg.scala 27:20]
  reg [63:0] _T_3_1_data; // @[Reg.scala 27:20]
  reg [63:0] _T_3_2_data; // @[Reg.scala 27:20]
  reg [63:0] _T_3_3_data; // @[Reg.scala 27:20]
  reg  _T_6; // @[SRAMTemplate.scala 130:58]
  reg [63:0] _T_8_0_data; // @[Reg.scala 27:20]
  reg [63:0] _T_8_1_data; // @[Reg.scala 27:20]
  reg [63:0] _T_8_2_data; // @[Reg.scala 27:20]
  reg [63:0] _T_8_3_data; // @[Reg.scala 27:20]
  SRAMTemplate_2 ram ( // @[SRAMTemplate.scala 121:19]
    .clock(ram_clock),
    .io_rreq_ready(ram_io_rreq_ready),
    .io_rreq_valid(ram_io_rreq_valid),
    .io_rreq_bits_setIdx(ram_io_rreq_bits_setIdx),
    .io_rresp_data_0_data(ram_io_rresp_data_0_data),
    .io_rresp_data_1_data(ram_io_rresp_data_1_data),
    .io_rresp_data_2_data(ram_io_rresp_data_2_data),
    .io_rresp_data_3_data(ram_io_rresp_data_3_data),
    .io_wreq_valid(ram_io_wreq_valid),
    .io_wreq_bits_setIdx(ram_io_wreq_bits_setIdx),
    .io_wreq_bits_data_data(ram_io_wreq_bits_data_data),
    .io_wreq_bits_waymask(ram_io_wreq_bits_waymask)
  );
  Arbiter_3 readArb ( // @[SRAMTemplate.scala 124:23]
    .io_in_0_ready(readArb_io_in_0_ready),
    .io_in_0_valid(readArb_io_in_0_valid),
    .io_in_0_bits_setIdx(readArb_io_in_0_bits_setIdx),
    .io_in_1_ready(readArb_io_in_1_ready),
    .io_in_1_valid(readArb_io_in_1_valid),
    .io_in_1_bits_setIdx(readArb_io_in_1_bits_setIdx),
    .io_out_ready(readArb_io_out_ready),
    .io_out_valid(readArb_io_out_valid),
    .io_out_bits_setIdx(readArb_io_out_bits_setIdx)
  );
  assign io_r0_req_ready = readArb_io_in_0_ready; // @[SRAMTemplate.scala 125:17]
  assign io_r0_resp_data_0_data = _T_1 ? ram_io_rresp_data_0_data : _T_3_0_data; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_1_data = _T_1 ? ram_io_rresp_data_1_data : _T_3_1_data; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_2_data = _T_1 ? ram_io_rresp_data_2_data : _T_3_2_data; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_3_data = _T_1 ? ram_io_rresp_data_3_data : _T_3_3_data; // @[SRAMTemplate.scala 130:17]
  assign io_r1_req_ready = readArb_io_in_1_ready; // @[SRAMTemplate.scala 125:17]
  assign io_r1_resp_data_0_data = _T_6 ? ram_io_rresp_data_0_data : _T_8_0_data; // @[SRAMTemplate.scala 130:17]
  assign io_r1_resp_data_1_data = _T_6 ? ram_io_rresp_data_1_data : _T_8_1_data; // @[SRAMTemplate.scala 130:17]
  assign io_r1_resp_data_2_data = _T_6 ? ram_io_rresp_data_2_data : _T_8_2_data; // @[SRAMTemplate.scala 130:17]
  assign io_r1_resp_data_3_data = _T_6 ? ram_io_rresp_data_3_data : _T_8_3_data; // @[SRAMTemplate.scala 130:17]
  assign ram_clock = clock;
  assign ram_io_rreq_valid = readArb_io_out_valid; // @[SRAMTemplate.scala 126:16]
  assign ram_io_rreq_bits_setIdx = readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 126:16]
  assign ram_io_wreq_valid = io_wreq_valid; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_setIdx = io_wreq_bits_setIdx; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_data_data = io_wreq_bits_data_data; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_waymask = io_wreq_bits_waymask; // @[SRAMTemplate.scala 122:12]
  assign readArb_io_in_0_valid = io_r0_req_valid; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_0_bits_setIdx = io_r0_req_bits_setIdx; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_1_valid = io_r1_req_valid; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_1_bits_setIdx = io_r1_req_bits_setIdx; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_out_ready = ram_io_rreq_ready; // @[SRAMTemplate.scala 126:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1 = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  _T_3_0_data = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  _T_3_1_data = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  _T_3_2_data = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  _T_3_3_data = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  _T_6 = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  _T_8_0_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  _T_8_1_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  _T_8_2_data = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  _T_8_3_data = _RAND_9[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_1 <= io_r0_req_ready & io_r0_req_valid;
    if (reset) begin
      _T_3_0_data <= 64'h0;
    end else if (_T_1) begin
      _T_3_0_data <= ram_io_rresp_data_0_data;
    end
    if (reset) begin
      _T_3_1_data <= 64'h0;
    end else if (_T_1) begin
      _T_3_1_data <= ram_io_rresp_data_1_data;
    end
    if (reset) begin
      _T_3_2_data <= 64'h0;
    end else if (_T_1) begin
      _T_3_2_data <= ram_io_rresp_data_2_data;
    end
    if (reset) begin
      _T_3_3_data <= 64'h0;
    end else if (_T_1) begin
      _T_3_3_data <= ram_io_rresp_data_3_data;
    end
    _T_6 <= io_r1_req_ready & io_r1_req_valid;
    if (reset) begin
      _T_8_0_data <= 64'h0;
    end else if (_T_6) begin
      _T_8_0_data <= ram_io_rresp_data_0_data;
    end
    if (reset) begin
      _T_8_1_data <= 64'h0;
    end else if (_T_6) begin
      _T_8_1_data <= ram_io_rresp_data_1_data;
    end
    if (reset) begin
      _T_8_2_data <= 64'h0;
    end else if (_T_6) begin
      _T_8_2_data <= ram_io_rresp_data_2_data;
    end
    if (reset) begin
      _T_8_3_data <= 64'h0;
    end else if (_T_6) begin
      _T_8_3_data <= ram_io_rresp_data_3_data;
    end
  end
endmodule
module Arbiter_4(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [86:0] io_in_0_bits_user,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [86:0] io_out_bits_user
);
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = io_in_0_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_addr = io_in_0_bits_addr; // @[Arbiter.scala 124:15]
  assign io_out_bits_user = io_in_0_bits_user; // @[Arbiter.scala 124:15]
endmodule
module Cache(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [86:0] io_in_req_bits_user,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  output [86:0] io_in_resp_bits_user,
  input  [1:0]  io_flush,
  input         io_out_mem_req_ready,
  output        io_out_mem_req_valid,
  output [31:0] io_out_mem_req_bits_addr,
  output [3:0]  io_out_mem_req_bits_cmd,
  output [63:0] io_out_mem_req_bits_wdata,
  input         io_out_mem_resp_valid,
  input  [3:0]  io_out_mem_resp_bits_cmd,
  input  [63:0] io_out_mem_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  input         io_mmio_resp_valid,
  input  [63:0] io_mmio_resp_bits_rdata,
  output        io_empty,
  input         MOUFlushICache
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [95:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [95:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [63:0] _RAND_18;
  reg [63:0] _RAND_19;
  reg [63:0] _RAND_20;
  reg [63:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [31:0] _RAND_27;
`endif // RANDOMIZE_REG_INIT
  wire  s1_io_in_ready; // @[Cache.scala 475:18]
  wire  s1_io_in_valid; // @[Cache.scala 475:18]
  wire [31:0] s1_io_in_bits_addr; // @[Cache.scala 475:18]
  wire [86:0] s1_io_in_bits_user; // @[Cache.scala 475:18]
  wire  s1_io_out_ready; // @[Cache.scala 475:18]
  wire  s1_io_out_valid; // @[Cache.scala 475:18]
  wire [31:0] s1_io_out_bits_req_addr; // @[Cache.scala 475:18]
  wire [86:0] s1_io_out_bits_req_user; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_req_ready; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_req_valid; // @[Cache.scala 475:18]
  wire [6:0] s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 475:18]
  wire [18:0] s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_0_dirty; // @[Cache.scala 475:18]
  wire [18:0] s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_1_dirty; // @[Cache.scala 475:18]
  wire [18:0] s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_2_dirty; // @[Cache.scala 475:18]
  wire [18:0] s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_3_dirty; // @[Cache.scala 475:18]
  wire  s1_io_dataReadBus_req_ready; // @[Cache.scala 475:18]
  wire  s1_io_dataReadBus_req_valid; // @[Cache.scala 475:18]
  wire [9:0] s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 475:18]
  wire [63:0] s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 475:18]
  wire [63:0] s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 475:18]
  wire [63:0] s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 475:18]
  wire [63:0] s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 475:18]
  wire  s2_clock; // @[Cache.scala 476:18]
  wire  s2_reset; // @[Cache.scala 476:18]
  wire  s2_io_in_ready; // @[Cache.scala 476:18]
  wire  s2_io_in_valid; // @[Cache.scala 476:18]
  wire [31:0] s2_io_in_bits_req_addr; // @[Cache.scala 476:18]
  wire [86:0] s2_io_in_bits_req_user; // @[Cache.scala 476:18]
  wire  s2_io_out_ready; // @[Cache.scala 476:18]
  wire  s2_io_out_valid; // @[Cache.scala 476:18]
  wire [31:0] s2_io_out_bits_req_addr; // @[Cache.scala 476:18]
  wire [86:0] s2_io_out_bits_req_user; // @[Cache.scala 476:18]
  wire [18:0] s2_io_out_bits_metas_0_tag; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_0_valid; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_0_dirty; // @[Cache.scala 476:18]
  wire [18:0] s2_io_out_bits_metas_1_tag; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_1_valid; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_1_dirty; // @[Cache.scala 476:18]
  wire [18:0] s2_io_out_bits_metas_2_tag; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_2_valid; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_2_dirty; // @[Cache.scala 476:18]
  wire [18:0] s2_io_out_bits_metas_3_tag; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_3_valid; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_3_dirty; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_datas_0_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_datas_1_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_datas_2_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_datas_3_data; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_hit; // @[Cache.scala 476:18]
  wire [3:0] s2_io_out_bits_waymask; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_mmio; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_isForwardData; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_forwardData_data_data; // @[Cache.scala 476:18]
  wire [3:0] s2_io_out_bits_forwardData_waymask; // @[Cache.scala 476:18]
  wire [18:0] s2_io_metaReadResp_0_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_0_valid; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_0_dirty; // @[Cache.scala 476:18]
  wire [18:0] s2_io_metaReadResp_1_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_1_valid; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_1_dirty; // @[Cache.scala 476:18]
  wire [18:0] s2_io_metaReadResp_2_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_2_valid; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_2_dirty; // @[Cache.scala 476:18]
  wire [18:0] s2_io_metaReadResp_3_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_3_valid; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_3_dirty; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataReadResp_0_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataReadResp_1_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataReadResp_2_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataReadResp_3_data; // @[Cache.scala 476:18]
  wire  s2_io_metaWriteBus_req_valid; // @[Cache.scala 476:18]
  wire [6:0] s2_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 476:18]
  wire [18:0] s2_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 476:18]
  wire [3:0] s2_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 476:18]
  wire  s2_io_dataWriteBus_req_valid; // @[Cache.scala 476:18]
  wire [9:0] s2_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 476:18]
  wire [3:0] s2_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 476:18]
  wire  s3_clock; // @[Cache.scala 477:18]
  wire  s3_reset; // @[Cache.scala 477:18]
  wire  s3_io_in_ready; // @[Cache.scala 477:18]
  wire  s3_io_in_valid; // @[Cache.scala 477:18]
  wire [31:0] s3_io_in_bits_req_addr; // @[Cache.scala 477:18]
  wire [86:0] s3_io_in_bits_req_user; // @[Cache.scala 477:18]
  wire [18:0] s3_io_in_bits_metas_0_tag; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_0_valid; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_0_dirty; // @[Cache.scala 477:18]
  wire [18:0] s3_io_in_bits_metas_1_tag; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_1_valid; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_1_dirty; // @[Cache.scala 477:18]
  wire [18:0] s3_io_in_bits_metas_2_tag; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_2_valid; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_2_dirty; // @[Cache.scala 477:18]
  wire [18:0] s3_io_in_bits_metas_3_tag; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_3_valid; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_3_dirty; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_datas_0_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_datas_1_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_datas_2_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_datas_3_data; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_hit; // @[Cache.scala 477:18]
  wire [3:0] s3_io_in_bits_waymask; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_mmio; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_isForwardData; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_forwardData_data_data; // @[Cache.scala 477:18]
  wire [3:0] s3_io_in_bits_forwardData_waymask; // @[Cache.scala 477:18]
  wire  s3_io_out_ready; // @[Cache.scala 477:18]
  wire  s3_io_out_valid; // @[Cache.scala 477:18]
  wire [63:0] s3_io_out_bits_rdata; // @[Cache.scala 477:18]
  wire [86:0] s3_io_out_bits_user; // @[Cache.scala 477:18]
  wire  s3_io_isFinish; // @[Cache.scala 477:18]
  wire  s3_io_flush; // @[Cache.scala 477:18]
  wire  s3_io_dataReadBus_req_ready; // @[Cache.scala 477:18]
  wire  s3_io_dataReadBus_req_valid; // @[Cache.scala 477:18]
  wire [9:0] s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataReadBus_resp_data_0_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataReadBus_resp_data_1_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataReadBus_resp_data_2_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataReadBus_resp_data_3_data; // @[Cache.scala 477:18]
  wire  s3_io_dataWriteBus_req_valid; // @[Cache.scala 477:18]
  wire [9:0] s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 477:18]
  wire [3:0] s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 477:18]
  wire  s3_io_metaWriteBus_req_valid; // @[Cache.scala 477:18]
  wire [6:0] s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 477:18]
  wire [18:0] s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 477:18]
  wire  s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 477:18]
  wire [3:0] s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 477:18]
  wire  s3_io_mem_req_ready; // @[Cache.scala 477:18]
  wire  s3_io_mem_req_valid; // @[Cache.scala 477:18]
  wire [31:0] s3_io_mem_req_bits_addr; // @[Cache.scala 477:18]
  wire [3:0] s3_io_mem_req_bits_cmd; // @[Cache.scala 477:18]
  wire [63:0] s3_io_mem_req_bits_wdata; // @[Cache.scala 477:18]
  wire  s3_io_mem_resp_ready; // @[Cache.scala 477:18]
  wire  s3_io_mem_resp_valid; // @[Cache.scala 477:18]
  wire [3:0] s3_io_mem_resp_bits_cmd; // @[Cache.scala 477:18]
  wire [63:0] s3_io_mem_resp_bits_rdata; // @[Cache.scala 477:18]
  wire  s3_io_mmio_req_ready; // @[Cache.scala 477:18]
  wire  s3_io_mmio_req_valid; // @[Cache.scala 477:18]
  wire [31:0] s3_io_mmio_req_bits_addr; // @[Cache.scala 477:18]
  wire  s3_io_mmio_resp_ready; // @[Cache.scala 477:18]
  wire  s3_io_mmio_resp_valid; // @[Cache.scala 477:18]
  wire [63:0] s3_io_mmio_resp_bits_rdata; // @[Cache.scala 477:18]
  wire  s3_io_cohResp_valid; // @[Cache.scala 477:18]
  wire  metaArray_clock; // @[Cache.scala 478:25]
  wire  metaArray_reset; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_req_ready; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_req_valid; // @[Cache.scala 478:25]
  wire [6:0] metaArray_io_r0_req_bits_setIdx; // @[Cache.scala 478:25]
  wire [18:0] metaArray_io_r0_resp_data_0_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_resp_data_0_valid; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_resp_data_0_dirty; // @[Cache.scala 478:25]
  wire [18:0] metaArray_io_r0_resp_data_1_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_resp_data_1_valid; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_resp_data_1_dirty; // @[Cache.scala 478:25]
  wire [18:0] metaArray_io_r0_resp_data_2_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_resp_data_2_valid; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_resp_data_2_dirty; // @[Cache.scala 478:25]
  wire [18:0] metaArray_io_r0_resp_data_3_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_resp_data_3_valid; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_resp_data_3_dirty; // @[Cache.scala 478:25]
  wire  metaArray_io_wreq_valid; // @[Cache.scala 478:25]
  wire [6:0] metaArray_io_wreq_bits_setIdx; // @[Cache.scala 478:25]
  wire [18:0] metaArray_io_wreq_bits_data_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_wreq_bits_data_dirty; // @[Cache.scala 478:25]
  wire [3:0] metaArray_io_wreq_bits_waymask; // @[Cache.scala 478:25]
  wire  dataArray_clock; // @[Cache.scala 479:25]
  wire  dataArray_reset; // @[Cache.scala 479:25]
  wire  dataArray_io_r0_req_ready; // @[Cache.scala 479:25]
  wire  dataArray_io_r0_req_valid; // @[Cache.scala 479:25]
  wire [9:0] dataArray_io_r0_req_bits_setIdx; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r0_resp_data_0_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r0_resp_data_1_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r0_resp_data_2_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r0_resp_data_3_data; // @[Cache.scala 479:25]
  wire  dataArray_io_r1_req_ready; // @[Cache.scala 479:25]
  wire  dataArray_io_r1_req_valid; // @[Cache.scala 479:25]
  wire [9:0] dataArray_io_r1_req_bits_setIdx; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r1_resp_data_0_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r1_resp_data_1_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r1_resp_data_2_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r1_resp_data_3_data; // @[Cache.scala 479:25]
  wire  dataArray_io_wreq_valid; // @[Cache.scala 479:25]
  wire [9:0] dataArray_io_wreq_bits_setIdx; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_wreq_bits_data_data; // @[Cache.scala 479:25]
  wire [3:0] dataArray_io_wreq_bits_waymask; // @[Cache.scala 479:25]
  wire  arb_io_in_0_ready; // @[Cache.scala 488:19]
  wire  arb_io_in_0_valid; // @[Cache.scala 488:19]
  wire [31:0] arb_io_in_0_bits_addr; // @[Cache.scala 488:19]
  wire [86:0] arb_io_in_0_bits_user; // @[Cache.scala 488:19]
  wire  arb_io_out_ready; // @[Cache.scala 488:19]
  wire  arb_io_out_valid; // @[Cache.scala 488:19]
  wire [31:0] arb_io_out_bits_addr; // @[Cache.scala 488:19]
  wire [86:0] arb_io_out_bits_user; // @[Cache.scala 488:19]
  wire  _T_3 = s2_io_out_ready & s2_io_out_valid; // @[Decoupled.scala 40:37]
  reg  _T_5; // @[Pipeline.scala 24:24]
  wire  _GEN_0 = _T_3 ? 1'h0 : _T_5; // @[Pipeline.scala 25:25]
  wire  _T_6 = s1_io_out_valid & s2_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_1 = _T_6 | _GEN_0; // @[Pipeline.scala 26:38]
  reg [31:0] _T_8_req_addr; // @[Reg.scala 15:16]
  reg [86:0] _T_8_req_user; // @[Reg.scala 15:16]
  reg  _T_10; // @[Pipeline.scala 24:24]
  wire  _GEN_9 = s3_io_isFinish ? 1'h0 : _T_10; // @[Pipeline.scala 25:25]
  wire  _T_11 = s2_io_out_valid & s3_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_10 = _T_11 | _GEN_9; // @[Pipeline.scala 26:38]
  reg [31:0] _T_13_req_addr; // @[Reg.scala 15:16]
  reg [86:0] _T_13_req_user; // @[Reg.scala 15:16]
  reg [18:0] _T_13_metas_0_tag; // @[Reg.scala 15:16]
  reg  _T_13_metas_0_valid; // @[Reg.scala 15:16]
  reg  _T_13_metas_0_dirty; // @[Reg.scala 15:16]
  reg [18:0] _T_13_metas_1_tag; // @[Reg.scala 15:16]
  reg  _T_13_metas_1_valid; // @[Reg.scala 15:16]
  reg  _T_13_metas_1_dirty; // @[Reg.scala 15:16]
  reg [18:0] _T_13_metas_2_tag; // @[Reg.scala 15:16]
  reg  _T_13_metas_2_valid; // @[Reg.scala 15:16]
  reg  _T_13_metas_2_dirty; // @[Reg.scala 15:16]
  reg [18:0] _T_13_metas_3_tag; // @[Reg.scala 15:16]
  reg  _T_13_metas_3_valid; // @[Reg.scala 15:16]
  reg  _T_13_metas_3_dirty; // @[Reg.scala 15:16]
  reg [63:0] _T_13_datas_0_data; // @[Reg.scala 15:16]
  reg [63:0] _T_13_datas_1_data; // @[Reg.scala 15:16]
  reg [63:0] _T_13_datas_2_data; // @[Reg.scala 15:16]
  reg [63:0] _T_13_datas_3_data; // @[Reg.scala 15:16]
  reg  _T_13_hit; // @[Reg.scala 15:16]
  reg [3:0] _T_13_waymask; // @[Reg.scala 15:16]
  reg  _T_13_mmio; // @[Reg.scala 15:16]
  reg  _T_13_isForwardData; // @[Reg.scala 15:16]
  reg [63:0] _T_13_forwardData_data_data; // @[Reg.scala 15:16]
  reg [3:0] _T_13_forwardData_waymask; // @[Reg.scala 15:16]
  wire  _T_15 = ~s2_io_in_valid; // @[Cache.scala 503:15]
  wire  _T_16 = ~s3_io_in_valid; // @[Cache.scala 503:34]
  CacheStage1 s1 ( // @[Cache.scala 475:18]
    .io_in_ready(s1_io_in_ready),
    .io_in_valid(s1_io_in_valid),
    .io_in_bits_addr(s1_io_in_bits_addr),
    .io_in_bits_user(s1_io_in_bits_user),
    .io_out_ready(s1_io_out_ready),
    .io_out_valid(s1_io_out_valid),
    .io_out_bits_req_addr(s1_io_out_bits_req_addr),
    .io_out_bits_req_user(s1_io_out_bits_req_user),
    .io_metaReadBus_req_ready(s1_io_metaReadBus_req_ready),
    .io_metaReadBus_req_valid(s1_io_metaReadBus_req_valid),
    .io_metaReadBus_req_bits_setIdx(s1_io_metaReadBus_req_bits_setIdx),
    .io_metaReadBus_resp_data_0_tag(s1_io_metaReadBus_resp_data_0_tag),
    .io_metaReadBus_resp_data_0_valid(s1_io_metaReadBus_resp_data_0_valid),
    .io_metaReadBus_resp_data_0_dirty(s1_io_metaReadBus_resp_data_0_dirty),
    .io_metaReadBus_resp_data_1_tag(s1_io_metaReadBus_resp_data_1_tag),
    .io_metaReadBus_resp_data_1_valid(s1_io_metaReadBus_resp_data_1_valid),
    .io_metaReadBus_resp_data_1_dirty(s1_io_metaReadBus_resp_data_1_dirty),
    .io_metaReadBus_resp_data_2_tag(s1_io_metaReadBus_resp_data_2_tag),
    .io_metaReadBus_resp_data_2_valid(s1_io_metaReadBus_resp_data_2_valid),
    .io_metaReadBus_resp_data_2_dirty(s1_io_metaReadBus_resp_data_2_dirty),
    .io_metaReadBus_resp_data_3_tag(s1_io_metaReadBus_resp_data_3_tag),
    .io_metaReadBus_resp_data_3_valid(s1_io_metaReadBus_resp_data_3_valid),
    .io_metaReadBus_resp_data_3_dirty(s1_io_metaReadBus_resp_data_3_dirty),
    .io_dataReadBus_req_ready(s1_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s1_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s1_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s1_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s1_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s1_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s1_io_dataReadBus_resp_data_3_data)
  );
  CacheStage2 s2 ( // @[Cache.scala 476:18]
    .clock(s2_clock),
    .reset(s2_reset),
    .io_in_ready(s2_io_in_ready),
    .io_in_valid(s2_io_in_valid),
    .io_in_bits_req_addr(s2_io_in_bits_req_addr),
    .io_in_bits_req_user(s2_io_in_bits_req_user),
    .io_out_ready(s2_io_out_ready),
    .io_out_valid(s2_io_out_valid),
    .io_out_bits_req_addr(s2_io_out_bits_req_addr),
    .io_out_bits_req_user(s2_io_out_bits_req_user),
    .io_out_bits_metas_0_tag(s2_io_out_bits_metas_0_tag),
    .io_out_bits_metas_0_valid(s2_io_out_bits_metas_0_valid),
    .io_out_bits_metas_0_dirty(s2_io_out_bits_metas_0_dirty),
    .io_out_bits_metas_1_tag(s2_io_out_bits_metas_1_tag),
    .io_out_bits_metas_1_valid(s2_io_out_bits_metas_1_valid),
    .io_out_bits_metas_1_dirty(s2_io_out_bits_metas_1_dirty),
    .io_out_bits_metas_2_tag(s2_io_out_bits_metas_2_tag),
    .io_out_bits_metas_2_valid(s2_io_out_bits_metas_2_valid),
    .io_out_bits_metas_2_dirty(s2_io_out_bits_metas_2_dirty),
    .io_out_bits_metas_3_tag(s2_io_out_bits_metas_3_tag),
    .io_out_bits_metas_3_valid(s2_io_out_bits_metas_3_valid),
    .io_out_bits_metas_3_dirty(s2_io_out_bits_metas_3_dirty),
    .io_out_bits_datas_0_data(s2_io_out_bits_datas_0_data),
    .io_out_bits_datas_1_data(s2_io_out_bits_datas_1_data),
    .io_out_bits_datas_2_data(s2_io_out_bits_datas_2_data),
    .io_out_bits_datas_3_data(s2_io_out_bits_datas_3_data),
    .io_out_bits_hit(s2_io_out_bits_hit),
    .io_out_bits_waymask(s2_io_out_bits_waymask),
    .io_out_bits_mmio(s2_io_out_bits_mmio),
    .io_out_bits_isForwardData(s2_io_out_bits_isForwardData),
    .io_out_bits_forwardData_data_data(s2_io_out_bits_forwardData_data_data),
    .io_out_bits_forwardData_waymask(s2_io_out_bits_forwardData_waymask),
    .io_metaReadResp_0_tag(s2_io_metaReadResp_0_tag),
    .io_metaReadResp_0_valid(s2_io_metaReadResp_0_valid),
    .io_metaReadResp_0_dirty(s2_io_metaReadResp_0_dirty),
    .io_metaReadResp_1_tag(s2_io_metaReadResp_1_tag),
    .io_metaReadResp_1_valid(s2_io_metaReadResp_1_valid),
    .io_metaReadResp_1_dirty(s2_io_metaReadResp_1_dirty),
    .io_metaReadResp_2_tag(s2_io_metaReadResp_2_tag),
    .io_metaReadResp_2_valid(s2_io_metaReadResp_2_valid),
    .io_metaReadResp_2_dirty(s2_io_metaReadResp_2_dirty),
    .io_metaReadResp_3_tag(s2_io_metaReadResp_3_tag),
    .io_metaReadResp_3_valid(s2_io_metaReadResp_3_valid),
    .io_metaReadResp_3_dirty(s2_io_metaReadResp_3_dirty),
    .io_dataReadResp_0_data(s2_io_dataReadResp_0_data),
    .io_dataReadResp_1_data(s2_io_dataReadResp_1_data),
    .io_dataReadResp_2_data(s2_io_dataReadResp_2_data),
    .io_dataReadResp_3_data(s2_io_dataReadResp_3_data),
    .io_metaWriteBus_req_valid(s2_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s2_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s2_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_dirty(s2_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s2_io_metaWriteBus_req_bits_waymask),
    .io_dataWriteBus_req_valid(s2_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s2_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s2_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s2_io_dataWriteBus_req_bits_waymask)
  );
  CacheStage3 s3 ( // @[Cache.scala 477:18]
    .clock(s3_clock),
    .reset(s3_reset),
    .io_in_ready(s3_io_in_ready),
    .io_in_valid(s3_io_in_valid),
    .io_in_bits_req_addr(s3_io_in_bits_req_addr),
    .io_in_bits_req_user(s3_io_in_bits_req_user),
    .io_in_bits_metas_0_tag(s3_io_in_bits_metas_0_tag),
    .io_in_bits_metas_0_valid(s3_io_in_bits_metas_0_valid),
    .io_in_bits_metas_0_dirty(s3_io_in_bits_metas_0_dirty),
    .io_in_bits_metas_1_tag(s3_io_in_bits_metas_1_tag),
    .io_in_bits_metas_1_valid(s3_io_in_bits_metas_1_valid),
    .io_in_bits_metas_1_dirty(s3_io_in_bits_metas_1_dirty),
    .io_in_bits_metas_2_tag(s3_io_in_bits_metas_2_tag),
    .io_in_bits_metas_2_valid(s3_io_in_bits_metas_2_valid),
    .io_in_bits_metas_2_dirty(s3_io_in_bits_metas_2_dirty),
    .io_in_bits_metas_3_tag(s3_io_in_bits_metas_3_tag),
    .io_in_bits_metas_3_valid(s3_io_in_bits_metas_3_valid),
    .io_in_bits_metas_3_dirty(s3_io_in_bits_metas_3_dirty),
    .io_in_bits_datas_0_data(s3_io_in_bits_datas_0_data),
    .io_in_bits_datas_1_data(s3_io_in_bits_datas_1_data),
    .io_in_bits_datas_2_data(s3_io_in_bits_datas_2_data),
    .io_in_bits_datas_3_data(s3_io_in_bits_datas_3_data),
    .io_in_bits_hit(s3_io_in_bits_hit),
    .io_in_bits_waymask(s3_io_in_bits_waymask),
    .io_in_bits_mmio(s3_io_in_bits_mmio),
    .io_in_bits_isForwardData(s3_io_in_bits_isForwardData),
    .io_in_bits_forwardData_data_data(s3_io_in_bits_forwardData_data_data),
    .io_in_bits_forwardData_waymask(s3_io_in_bits_forwardData_waymask),
    .io_out_ready(s3_io_out_ready),
    .io_out_valid(s3_io_out_valid),
    .io_out_bits_rdata(s3_io_out_bits_rdata),
    .io_out_bits_user(s3_io_out_bits_user),
    .io_isFinish(s3_io_isFinish),
    .io_flush(s3_io_flush),
    .io_dataReadBus_req_ready(s3_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s3_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s3_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s3_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s3_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s3_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s3_io_dataReadBus_resp_data_3_data),
    .io_dataWriteBus_req_valid(s3_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s3_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s3_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s3_io_dataWriteBus_req_bits_waymask),
    .io_metaWriteBus_req_valid(s3_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s3_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s3_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_dirty(s3_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s3_io_metaWriteBus_req_bits_waymask),
    .io_mem_req_ready(s3_io_mem_req_ready),
    .io_mem_req_valid(s3_io_mem_req_valid),
    .io_mem_req_bits_addr(s3_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(s3_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(s3_io_mem_req_bits_wdata),
    .io_mem_resp_ready(s3_io_mem_resp_ready),
    .io_mem_resp_valid(s3_io_mem_resp_valid),
    .io_mem_resp_bits_cmd(s3_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_rdata(s3_io_mem_resp_bits_rdata),
    .io_mmio_req_ready(s3_io_mmio_req_ready),
    .io_mmio_req_valid(s3_io_mmio_req_valid),
    .io_mmio_req_bits_addr(s3_io_mmio_req_bits_addr),
    .io_mmio_resp_ready(s3_io_mmio_resp_ready),
    .io_mmio_resp_valid(s3_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(s3_io_mmio_resp_bits_rdata),
    .io_cohResp_valid(s3_io_cohResp_valid)
  );
  SRAMTemplateWithArbiter metaArray ( // @[Cache.scala 478:25]
    .clock(metaArray_clock),
    .reset(metaArray_reset),
    .io_r0_req_ready(metaArray_io_r0_req_ready),
    .io_r0_req_valid(metaArray_io_r0_req_valid),
    .io_r0_req_bits_setIdx(metaArray_io_r0_req_bits_setIdx),
    .io_r0_resp_data_0_tag(metaArray_io_r0_resp_data_0_tag),
    .io_r0_resp_data_0_valid(metaArray_io_r0_resp_data_0_valid),
    .io_r0_resp_data_0_dirty(metaArray_io_r0_resp_data_0_dirty),
    .io_r0_resp_data_1_tag(metaArray_io_r0_resp_data_1_tag),
    .io_r0_resp_data_1_valid(metaArray_io_r0_resp_data_1_valid),
    .io_r0_resp_data_1_dirty(metaArray_io_r0_resp_data_1_dirty),
    .io_r0_resp_data_2_tag(metaArray_io_r0_resp_data_2_tag),
    .io_r0_resp_data_2_valid(metaArray_io_r0_resp_data_2_valid),
    .io_r0_resp_data_2_dirty(metaArray_io_r0_resp_data_2_dirty),
    .io_r0_resp_data_3_tag(metaArray_io_r0_resp_data_3_tag),
    .io_r0_resp_data_3_valid(metaArray_io_r0_resp_data_3_valid),
    .io_r0_resp_data_3_dirty(metaArray_io_r0_resp_data_3_dirty),
    .io_wreq_valid(metaArray_io_wreq_valid),
    .io_wreq_bits_setIdx(metaArray_io_wreq_bits_setIdx),
    .io_wreq_bits_data_tag(metaArray_io_wreq_bits_data_tag),
    .io_wreq_bits_data_dirty(metaArray_io_wreq_bits_data_dirty),
    .io_wreq_bits_waymask(metaArray_io_wreq_bits_waymask)
  );
  SRAMTemplateWithArbiter_1 dataArray ( // @[Cache.scala 479:25]
    .clock(dataArray_clock),
    .reset(dataArray_reset),
    .io_r0_req_ready(dataArray_io_r0_req_ready),
    .io_r0_req_valid(dataArray_io_r0_req_valid),
    .io_r0_req_bits_setIdx(dataArray_io_r0_req_bits_setIdx),
    .io_r0_resp_data_0_data(dataArray_io_r0_resp_data_0_data),
    .io_r0_resp_data_1_data(dataArray_io_r0_resp_data_1_data),
    .io_r0_resp_data_2_data(dataArray_io_r0_resp_data_2_data),
    .io_r0_resp_data_3_data(dataArray_io_r0_resp_data_3_data),
    .io_r1_req_ready(dataArray_io_r1_req_ready),
    .io_r1_req_valid(dataArray_io_r1_req_valid),
    .io_r1_req_bits_setIdx(dataArray_io_r1_req_bits_setIdx),
    .io_r1_resp_data_0_data(dataArray_io_r1_resp_data_0_data),
    .io_r1_resp_data_1_data(dataArray_io_r1_resp_data_1_data),
    .io_r1_resp_data_2_data(dataArray_io_r1_resp_data_2_data),
    .io_r1_resp_data_3_data(dataArray_io_r1_resp_data_3_data),
    .io_wreq_valid(dataArray_io_wreq_valid),
    .io_wreq_bits_setIdx(dataArray_io_wreq_bits_setIdx),
    .io_wreq_bits_data_data(dataArray_io_wreq_bits_data_data),
    .io_wreq_bits_waymask(dataArray_io_wreq_bits_waymask)
  );
  Arbiter_4 arb ( // @[Cache.scala 488:19]
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_addr(arb_io_in_0_bits_addr),
    .io_in_0_bits_user(arb_io_in_0_bits_user),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_addr(arb_io_out_bits_addr),
    .io_out_bits_user(arb_io_out_bits_user)
  );
  assign io_in_req_ready = arb_io_in_0_ready; // @[Cache.scala 489:28]
  assign io_in_resp_valid = s3_io_out_valid; // @[Cache.scala 499:14 Cache.scala 505:20]
  assign io_in_resp_bits_rdata = s3_io_out_bits_rdata; // @[Cache.scala 499:14]
  assign io_in_resp_bits_user = s3_io_out_bits_user; // @[Cache.scala 499:14]
  assign io_out_mem_req_valid = s3_io_mem_req_valid; // @[Cache.scala 501:14]
  assign io_out_mem_req_bits_addr = s3_io_mem_req_bits_addr; // @[Cache.scala 501:14]
  assign io_out_mem_req_bits_cmd = s3_io_mem_req_bits_cmd; // @[Cache.scala 501:14]
  assign io_out_mem_req_bits_wdata = s3_io_mem_req_bits_wdata; // @[Cache.scala 501:14]
  assign io_mmio_req_valid = s3_io_mmio_req_valid; // @[Cache.scala 502:11]
  assign io_mmio_req_bits_addr = s3_io_mmio_req_bits_addr; // @[Cache.scala 502:11]
  assign io_empty = _T_15 & _T_16; // @[Cache.scala 503:12]
  assign s1_io_in_valid = arb_io_out_valid; // @[Cache.scala 491:12]
  assign s1_io_in_bits_addr = arb_io_out_bits_addr; // @[Cache.scala 491:12]
  assign s1_io_in_bits_user = arb_io_out_bits_user; // @[Cache.scala 491:12]
  assign s1_io_out_ready = s2_io_in_ready; // @[Pipeline.scala 29:16]
  assign s1_io_metaReadBus_req_ready = metaArray_io_r0_req_ready; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_0_tag = metaArray_io_r0_resp_data_0_tag; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_0_valid = metaArray_io_r0_resp_data_0_valid; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_0_dirty = metaArray_io_r0_resp_data_0_dirty; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_1_tag = metaArray_io_r0_resp_data_1_tag; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_1_valid = metaArray_io_r0_resp_data_1_valid; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_1_dirty = metaArray_io_r0_resp_data_1_dirty; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_2_tag = metaArray_io_r0_resp_data_2_tag; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_2_valid = metaArray_io_r0_resp_data_2_valid; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_2_dirty = metaArray_io_r0_resp_data_2_dirty; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_3_tag = metaArray_io_r0_resp_data_3_tag; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_3_valid = metaArray_io_r0_resp_data_3_valid; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_3_dirty = metaArray_io_r0_resp_data_3_dirty; // @[Cache.scala 523:21]
  assign s1_io_dataReadBus_req_ready = dataArray_io_r0_req_ready; // @[Cache.scala 524:21]
  assign s1_io_dataReadBus_resp_data_0_data = dataArray_io_r0_resp_data_0_data; // @[Cache.scala 524:21]
  assign s1_io_dataReadBus_resp_data_1_data = dataArray_io_r0_resp_data_1_data; // @[Cache.scala 524:21]
  assign s1_io_dataReadBus_resp_data_2_data = dataArray_io_r0_resp_data_2_data; // @[Cache.scala 524:21]
  assign s1_io_dataReadBus_resp_data_3_data = dataArray_io_r0_resp_data_3_data; // @[Cache.scala 524:21]
  assign s2_clock = clock;
  assign s2_reset = reset;
  assign s2_io_in_valid = _T_5; // @[Pipeline.scala 31:17]
  assign s2_io_in_bits_req_addr = _T_8_req_addr; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_user = _T_8_req_user; // @[Pipeline.scala 30:16]
  assign s2_io_out_ready = s3_io_in_ready; // @[Pipeline.scala 29:16]
  assign s2_io_metaReadResp_0_tag = s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_0_valid = s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_0_dirty = s1_io_metaReadBus_resp_data_0_dirty; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_1_tag = s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_1_valid = s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_1_dirty = s1_io_metaReadBus_resp_data_1_dirty; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_2_tag = s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_2_valid = s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_2_dirty = s1_io_metaReadBus_resp_data_2_dirty; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_3_tag = s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_3_valid = s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_3_dirty = s1_io_metaReadBus_resp_data_3_dirty; // @[Cache.scala 530:22]
  assign s2_io_dataReadResp_0_data = s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 531:22]
  assign s2_io_dataReadResp_1_data = s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 531:22]
  assign s2_io_dataReadResp_2_data = s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 531:22]
  assign s2_io_dataReadResp_3_data = s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 531:22]
  assign s2_io_metaWriteBus_req_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 533:22]
  assign s2_io_metaWriteBus_req_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 533:22]
  assign s2_io_metaWriteBus_req_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 533:22]
  assign s2_io_metaWriteBus_req_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 533:22]
  assign s2_io_metaWriteBus_req_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 533:22]
  assign s2_io_dataWriteBus_req_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 532:22]
  assign s2_io_dataWriteBus_req_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 532:22]
  assign s2_io_dataWriteBus_req_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 532:22]
  assign s2_io_dataWriteBus_req_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 532:22]
  assign s3_clock = clock;
  assign s3_reset = reset;
  assign s3_io_in_valid = _T_10; // @[Pipeline.scala 31:17]
  assign s3_io_in_bits_req_addr = _T_13_req_addr; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_user = _T_13_req_user; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_tag = _T_13_metas_0_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_valid = _T_13_metas_0_valid; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_dirty = _T_13_metas_0_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_tag = _T_13_metas_1_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_valid = _T_13_metas_1_valid; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_dirty = _T_13_metas_1_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_tag = _T_13_metas_2_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_valid = _T_13_metas_2_valid; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_dirty = _T_13_metas_2_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_tag = _T_13_metas_3_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_valid = _T_13_metas_3_valid; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_dirty = _T_13_metas_3_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_0_data = _T_13_datas_0_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_1_data = _T_13_datas_1_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_2_data = _T_13_datas_2_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_3_data = _T_13_datas_3_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_hit = _T_13_hit; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_waymask = _T_13_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_mmio = _T_13_mmio; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_isForwardData = _T_13_isForwardData; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_data_data = _T_13_forwardData_data_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_waymask = _T_13_forwardData_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_out_ready = io_in_resp_ready; // @[Cache.scala 499:14]
  assign s3_io_flush = io_flush[1]; // @[Cache.scala 500:15]
  assign s3_io_dataReadBus_req_ready = dataArray_io_r1_req_ready; // @[Cache.scala 525:21]
  assign s3_io_dataReadBus_resp_data_0_data = dataArray_io_r1_resp_data_0_data; // @[Cache.scala 525:21]
  assign s3_io_dataReadBus_resp_data_1_data = dataArray_io_r1_resp_data_1_data; // @[Cache.scala 525:21]
  assign s3_io_dataReadBus_resp_data_2_data = dataArray_io_r1_resp_data_2_data; // @[Cache.scala 525:21]
  assign s3_io_dataReadBus_resp_data_3_data = dataArray_io_r1_resp_data_3_data; // @[Cache.scala 525:21]
  assign s3_io_mem_req_ready = io_out_mem_req_ready; // @[Cache.scala 501:14]
  assign s3_io_mem_resp_valid = io_out_mem_resp_valid; // @[Cache.scala 501:14]
  assign s3_io_mem_resp_bits_cmd = io_out_mem_resp_bits_cmd; // @[Cache.scala 501:14]
  assign s3_io_mem_resp_bits_rdata = io_out_mem_resp_bits_rdata; // @[Cache.scala 501:14]
  assign s3_io_mmio_req_ready = io_mmio_req_ready; // @[Cache.scala 502:11]
  assign s3_io_mmio_resp_valid = io_mmio_resp_valid; // @[Cache.scala 502:11]
  assign s3_io_mmio_resp_bits_rdata = io_mmio_resp_bits_rdata; // @[Cache.scala 502:11]
  assign metaArray_clock = clock;
  assign metaArray_reset = reset | MOUFlushICache; // @[Cache.scala 485:21]
  assign metaArray_io_r0_req_valid = s1_io_metaReadBus_req_valid; // @[Cache.scala 523:21]
  assign metaArray_io_r0_req_bits_setIdx = s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 523:21]
  assign metaArray_io_wreq_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 527:18]
  assign metaArray_io_wreq_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 527:18]
  assign metaArray_io_wreq_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 527:18]
  assign metaArray_io_wreq_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 527:18]
  assign metaArray_io_wreq_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 527:18]
  assign dataArray_clock = clock;
  assign dataArray_reset = reset;
  assign dataArray_io_r0_req_valid = s1_io_dataReadBus_req_valid; // @[Cache.scala 524:21]
  assign dataArray_io_r0_req_bits_setIdx = s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 524:21]
  assign dataArray_io_r1_req_valid = s3_io_dataReadBus_req_valid; // @[Cache.scala 525:21]
  assign dataArray_io_r1_req_bits_setIdx = s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 525:21]
  assign dataArray_io_wreq_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 528:18]
  assign dataArray_io_wreq_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 528:18]
  assign dataArray_io_wreq_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 528:18]
  assign dataArray_io_wreq_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 528:18]
  assign arb_io_in_0_valid = io_in_req_valid; // @[Cache.scala 489:28]
  assign arb_io_in_0_bits_addr = io_in_req_bits_addr; // @[Cache.scala 489:28]
  assign arb_io_in_0_bits_user = io_in_req_bits_user; // @[Cache.scala 489:28]
  assign arb_io_out_ready = s1_io_in_ready; // @[Cache.scala 491:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_5 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _T_8_req_addr = _RAND_1[31:0];
  _RAND_2 = {3{`RANDOM}};
  _T_8_req_user = _RAND_2[86:0];
  _RAND_3 = {1{`RANDOM}};
  _T_10 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_13_req_addr = _RAND_4[31:0];
  _RAND_5 = {3{`RANDOM}};
  _T_13_req_user = _RAND_5[86:0];
  _RAND_6 = {1{`RANDOM}};
  _T_13_metas_0_tag = _RAND_6[18:0];
  _RAND_7 = {1{`RANDOM}};
  _T_13_metas_0_valid = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_13_metas_0_dirty = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _T_13_metas_1_tag = _RAND_9[18:0];
  _RAND_10 = {1{`RANDOM}};
  _T_13_metas_1_valid = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_13_metas_1_dirty = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _T_13_metas_2_tag = _RAND_12[18:0];
  _RAND_13 = {1{`RANDOM}};
  _T_13_metas_2_valid = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _T_13_metas_2_dirty = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _T_13_metas_3_tag = _RAND_15[18:0];
  _RAND_16 = {1{`RANDOM}};
  _T_13_metas_3_valid = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  _T_13_metas_3_dirty = _RAND_17[0:0];
  _RAND_18 = {2{`RANDOM}};
  _T_13_datas_0_data = _RAND_18[63:0];
  _RAND_19 = {2{`RANDOM}};
  _T_13_datas_1_data = _RAND_19[63:0];
  _RAND_20 = {2{`RANDOM}};
  _T_13_datas_2_data = _RAND_20[63:0];
  _RAND_21 = {2{`RANDOM}};
  _T_13_datas_3_data = _RAND_21[63:0];
  _RAND_22 = {1{`RANDOM}};
  _T_13_hit = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  _T_13_waymask = _RAND_23[3:0];
  _RAND_24 = {1{`RANDOM}};
  _T_13_mmio = _RAND_24[0:0];
  _RAND_25 = {1{`RANDOM}};
  _T_13_isForwardData = _RAND_25[0:0];
  _RAND_26 = {2{`RANDOM}};
  _T_13_forwardData_data_data = _RAND_26[63:0];
  _RAND_27 = {1{`RANDOM}};
  _T_13_forwardData_waymask = _RAND_27[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_5 <= 1'h0;
    end else if (io_flush[0]) begin
      _T_5 <= 1'h0;
    end else begin
      _T_5 <= _GEN_1;
    end
    if (_T_6) begin
      _T_8_req_addr <= s1_io_out_bits_req_addr;
    end
    if (_T_6) begin
      _T_8_req_user <= s1_io_out_bits_req_user;
    end
    if (reset) begin
      _T_10 <= 1'h0;
    end else if (io_flush[1]) begin
      _T_10 <= 1'h0;
    end else begin
      _T_10 <= _GEN_10;
    end
    if (_T_11) begin
      _T_13_req_addr <= s2_io_out_bits_req_addr;
    end
    if (_T_11) begin
      _T_13_req_user <= s2_io_out_bits_req_user;
    end
    if (_T_11) begin
      _T_13_metas_0_tag <= s2_io_out_bits_metas_0_tag;
    end
    if (_T_11) begin
      _T_13_metas_0_valid <= s2_io_out_bits_metas_0_valid;
    end
    if (_T_11) begin
      _T_13_metas_0_dirty <= s2_io_out_bits_metas_0_dirty;
    end
    if (_T_11) begin
      _T_13_metas_1_tag <= s2_io_out_bits_metas_1_tag;
    end
    if (_T_11) begin
      _T_13_metas_1_valid <= s2_io_out_bits_metas_1_valid;
    end
    if (_T_11) begin
      _T_13_metas_1_dirty <= s2_io_out_bits_metas_1_dirty;
    end
    if (_T_11) begin
      _T_13_metas_2_tag <= s2_io_out_bits_metas_2_tag;
    end
    if (_T_11) begin
      _T_13_metas_2_valid <= s2_io_out_bits_metas_2_valid;
    end
    if (_T_11) begin
      _T_13_metas_2_dirty <= s2_io_out_bits_metas_2_dirty;
    end
    if (_T_11) begin
      _T_13_metas_3_tag <= s2_io_out_bits_metas_3_tag;
    end
    if (_T_11) begin
      _T_13_metas_3_valid <= s2_io_out_bits_metas_3_valid;
    end
    if (_T_11) begin
      _T_13_metas_3_dirty <= s2_io_out_bits_metas_3_dirty;
    end
    if (_T_11) begin
      _T_13_datas_0_data <= s2_io_out_bits_datas_0_data;
    end
    if (_T_11) begin
      _T_13_datas_1_data <= s2_io_out_bits_datas_1_data;
    end
    if (_T_11) begin
      _T_13_datas_2_data <= s2_io_out_bits_datas_2_data;
    end
    if (_T_11) begin
      _T_13_datas_3_data <= s2_io_out_bits_datas_3_data;
    end
    if (_T_11) begin
      _T_13_hit <= s2_io_out_bits_hit;
    end
    if (_T_11) begin
      _T_13_waymask <= s2_io_out_bits_waymask;
    end
    if (_T_11) begin
      _T_13_mmio <= s2_io_out_bits_mmio;
    end
    if (_T_11) begin
      _T_13_isForwardData <= s2_io_out_bits_isForwardData;
    end
    if (_T_11) begin
      _T_13_forwardData_data_data <= s2_io_out_bits_forwardData_data_data;
    end
    if (_T_11) begin
      _T_13_forwardData_waymask <= s2_io_out_bits_forwardData_waymask;
    end
  end
endmodule
module EmbeddedTLBExec_1(
  input          clock,
  input          reset,
  output         io_in_ready,
  input          io_in_valid,
  input  [38:0]  io_in_bits_addr,
  input  [2:0]   io_in_bits_size,
  input  [3:0]   io_in_bits_cmd,
  input  [7:0]   io_in_bits_wmask,
  input  [63:0]  io_in_bits_wdata,
  input          io_out_ready,
  output         io_out_valid,
  output [31:0]  io_out_bits_addr,
  output [2:0]   io_out_bits_size,
  output [3:0]   io_out_bits_cmd,
  output [7:0]   io_out_bits_wmask,
  output [63:0]  io_out_bits_wdata,
  input  [120:0] io_md_0,
  input  [120:0] io_md_1,
  input  [120:0] io_md_2,
  input  [120:0] io_md_3,
  output         io_mdWrite_wen,
  output [3:0]   io_mdWrite_windex,
  output [3:0]   io_mdWrite_waymask,
  output [120:0] io_mdWrite_wdata,
  input          io_mdReady,
  input          io_mem_req_ready,
  output         io_mem_req_valid,
  output [31:0]  io_mem_req_bits_addr,
  output [3:0]   io_mem_req_bits_cmd,
  output [63:0]  io_mem_req_bits_wdata,
  output         io_mem_resp_ready,
  input          io_mem_resp_valid,
  input  [63:0]  io_mem_resp_bits_rdata,
  input  [63:0]  io_satp,
  input  [1:0]   io_pf_priviledgeMode,
  input          io_pf_status_sum,
  input          io_pf_status_mxr,
  output         io_pf_loadPF,
  output         io_pf_storePF,
  output [38:0]  io_pf_addr,
  output         io_isFinish,
  input          ISAMO
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
`endif // RANDOMIZE_REG_INIT
  wire [8:0] vpn_vpn0 = io_in_bits_addr[20:12]; // @[EmbeddedTLB.scala 193:54]
  wire [8:0] vpn_vpn1 = io_in_bits_addr[29:21]; // @[EmbeddedTLB.scala 193:54]
  wire [8:0] vpn_vpn2 = io_in_bits_addr[38:30]; // @[EmbeddedTLB.scala 193:54]
  wire [19:0] satp_ppn = io_satp[19:0]; // @[EmbeddedTLB.scala 195:30]
  wire [15:0] satp_asid = io_satp[59:44]; // @[EmbeddedTLB.scala 195:30]
  wire  _T_39 = io_md_0[93:78] == satp_asid; // @[EmbeddedTLB.scala 204:117]
  wire  _T_40 = io_md_0[52] & _T_39; // @[EmbeddedTLB.scala 204:86]
  wire [17:0] _T_57 = {vpn_vpn2,vpn_vpn1}; // @[EmbeddedTLB.scala 204:201]
  wire [26:0] _T_58 = {vpn_vpn2,vpn_vpn1,vpn_vpn0}; // @[EmbeddedTLB.scala 204:201]
  wire [26:0] _T_59 = {9'h1ff,io_md_0[77:60]}; // @[Cat.scala 29:58]
  wire [26:0] _T_60 = _T_59 & io_md_0[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_62 = _T_59 & _T_58; // @[TLB.scala 131:84]
  wire  _T_63 = _T_60 == _T_62; // @[TLB.scala 131:48]
  wire  _T_64 = _T_40 & _T_63; // @[EmbeddedTLB.scala 204:132]
  wire  _T_91 = io_md_1[93:78] == satp_asid; // @[EmbeddedTLB.scala 204:117]
  wire  _T_92 = io_md_1[52] & _T_91; // @[EmbeddedTLB.scala 204:86]
  wire [26:0] _T_111 = {9'h1ff,io_md_1[77:60]}; // @[Cat.scala 29:58]
  wire [26:0] _T_112 = _T_111 & io_md_1[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_114 = _T_111 & _T_58; // @[TLB.scala 131:84]
  wire  _T_115 = _T_112 == _T_114; // @[TLB.scala 131:48]
  wire  _T_116 = _T_92 & _T_115; // @[EmbeddedTLB.scala 204:132]
  wire  _T_143 = io_md_2[93:78] == satp_asid; // @[EmbeddedTLB.scala 204:117]
  wire  _T_144 = io_md_2[52] & _T_143; // @[EmbeddedTLB.scala 204:86]
  wire [26:0] _T_163 = {9'h1ff,io_md_2[77:60]}; // @[Cat.scala 29:58]
  wire [26:0] _T_164 = _T_163 & io_md_2[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_166 = _T_163 & _T_58; // @[TLB.scala 131:84]
  wire  _T_167 = _T_164 == _T_166; // @[TLB.scala 131:48]
  wire  _T_168 = _T_144 & _T_167; // @[EmbeddedTLB.scala 204:132]
  wire  _T_195 = io_md_3[93:78] == satp_asid; // @[EmbeddedTLB.scala 204:117]
  wire  _T_196 = io_md_3[52] & _T_195; // @[EmbeddedTLB.scala 204:86]
  wire [26:0] _T_215 = {9'h1ff,io_md_3[77:60]}; // @[Cat.scala 29:58]
  wire [26:0] _T_216 = _T_215 & io_md_3[120:94]; // @[TLB.scala 131:37]
  wire [26:0] _T_218 = _T_215 & _T_58; // @[TLB.scala 131:84]
  wire  _T_219 = _T_216 == _T_218; // @[TLB.scala 131:48]
  wire  _T_220 = _T_196 & _T_219; // @[EmbeddedTLB.scala 204:132]
  wire [3:0] hitVec = {_T_220,_T_168,_T_116,_T_64}; // @[EmbeddedTLB.scala 204:211]
  wire  _T_224 = |hitVec; // @[EmbeddedTLB.scala 205:35]
  wire  hit = io_in_valid & _T_224; // @[EmbeddedTLB.scala 205:25]
  wire  _T_226 = ~_T_224; // @[EmbeddedTLB.scala 206:29]
  wire  miss = io_in_valid & _T_226; // @[EmbeddedTLB.scala 206:26]
  reg [63:0] _T_227; // @[LFSR64.scala 25:23]
  wire  _T_230 = _T_227[0] ^ _T_227[1]; // @[LFSR64.scala 26:23]
  wire  _T_232 = _T_230 ^ _T_227[3]; // @[LFSR64.scala 26:33]
  wire  _T_234 = _T_232 ^ _T_227[4]; // @[LFSR64.scala 26:43]
  wire  _T_235 = _T_227 == 64'h0; // @[LFSR64.scala 28:24]
  wire [63:0] _T_237 = {_T_234,_T_227[63:1]}; // @[Cat.scala 29:58]
  wire [3:0] victimWaymask = 4'h1 << _T_227[1:0]; // @[EmbeddedTLB.scala 208:42]
  wire [3:0] waymask = hit ? hitVec : victimWaymask; // @[EmbeddedTLB.scala 209:20]
  wire [120:0] _T_244 = waymask[0] ? io_md_0 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_245 = waymask[1] ? io_md_1 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_246 = waymask[2] ? io_md_2 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_247 = waymask[3] ? io_md_3 : 121'h0; // @[Mux.scala 27:72]
  wire [120:0] _T_248 = _T_244 | _T_245; // @[Mux.scala 27:72]
  wire [120:0] _T_249 = _T_248 | _T_246; // @[Mux.scala 27:72]
  wire [120:0] _T_250 = _T_249 | _T_247; // @[Mux.scala 27:72]
  wire [7:0] hitMeta_flag = _T_250[59:52]; // @[EmbeddedTLB.scala 215:70]
  wire [17:0] hitMeta_mask = _T_250[77:60]; // @[EmbeddedTLB.scala 215:70]
  wire [15:0] hitMeta_asid = _T_250[93:78]; // @[EmbeddedTLB.scala 215:70]
  wire [31:0] hitData_pteaddr = _T_250[31:0]; // @[EmbeddedTLB.scala 216:70]
  wire [19:0] hitData_ppn = _T_250[51:32]; // @[EmbeddedTLB.scala 216:70]
  wire  hitFlag_v = hitMeta_flag[0]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_r = hitMeta_flag[1]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_w = hitMeta_flag[2]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_x = hitMeta_flag[3]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_u = hitMeta_flag[4]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_g = hitMeta_flag[5]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_a = hitMeta_flag[6]; // @[EmbeddedTLB.scala 217:38]
  wire  hitFlag_d = hitMeta_flag[7]; // @[EmbeddedTLB.scala 217:38]
  wire  _T_289 = ~hitFlag_a; // @[EmbeddedTLB.scala 221:23]
  wire  _T_290 = ~hitFlag_d; // @[EmbeddedTLB.scala 221:37]
  wire  _T_292 = _T_290 & io_in_bits_cmd[0]; // @[EmbeddedTLB.scala 221:48]
  wire  _T_293 = _T_289 | _T_292; // @[EmbeddedTLB.scala 221:34]
  wire  _T_294 = hit & _T_293; // @[EmbeddedTLB.scala 221:19]
  reg [2:0] state; // @[EmbeddedTLB.scala 247:22]
  wire  _T_370 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_314 = io_pf_priviledgeMode == 2'h0; // @[EmbeddedTLB.scala 226:62]
  wire  _T_315 = ~hitFlag_u; // @[EmbeddedTLB.scala 226:75]
  wire  _T_316 = _T_314 & _T_315; // @[EmbeddedTLB.scala 226:72]
  wire  _T_317 = ~_T_316; // @[EmbeddedTLB.scala 226:42]
  wire  _T_318 = hit & _T_317; // @[EmbeddedTLB.scala 226:39]
  wire  _T_319 = io_pf_priviledgeMode == 2'h1; // @[EmbeddedTLB.scala 226:110]
  wire  _T_320 = _T_319 & hitFlag_u; // @[EmbeddedTLB.scala 226:120]
  wire  _T_321 = ~io_pf_status_sum; // @[EmbeddedTLB.scala 226:137]
  wire  _T_323 = _T_320 & _T_321; // @[EmbeddedTLB.scala 226:133]
  wire  _T_324 = ~_T_323; // @[EmbeddedTLB.scala 226:90]
  wire  hitCheck = _T_318 & _T_324; // @[EmbeddedTLB.scala 226:87]
  wire  _T_325 = io_pf_status_mxr & hitFlag_x; // @[EmbeddedTLB.scala 228:57]
  wire  _T_326 = hitFlag_r | _T_325; // @[EmbeddedTLB.scala 228:40]
  wire  hitLoad = hitCheck & _T_326; // @[EmbeddedTLB.scala 228:26]
  wire  _T_329 = ~hitLoad; // @[EmbeddedTLB.scala 241:15]
  wire  _T_331 = ~io_in_bits_cmd[0]; // @[SimpleBus.scala 73:18]
  wire  _T_333 = ~io_in_bits_cmd[3]; // @[SimpleBus.scala 73:29]
  wire  _T_334 = _T_331 & _T_333; // @[SimpleBus.scala 73:26]
  wire  _T_335 = _T_329 & _T_334; // @[EmbeddedTLB.scala 241:24]
  wire  _T_336 = _T_335 & hit; // @[EmbeddedTLB.scala 241:40]
  wire  _T_337 = ~ISAMO; // @[EmbeddedTLB.scala 241:50]
  wire  _T_338 = _T_336 & _T_337; // @[EmbeddedTLB.scala 241:47]
  wire  _T_377 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_379 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_397 = io_mem_resp_ready & io_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  memRdata_flag_d = io_mem_resp_bits_rdata[7]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_a = io_mem_resp_bits_rdata[6]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_g = io_mem_resp_bits_rdata[5]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_u = io_mem_resp_bits_rdata[4]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_x = io_mem_resp_bits_rdata[3]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_w = io_mem_resp_bits_rdata[2]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_r = io_mem_resp_bits_rdata[1]; // @[EmbeddedTLB.scala 255:49]
  wire  memRdata_flag_v = io_mem_resp_bits_rdata[0]; // @[EmbeddedTLB.scala 255:49]
  wire [7:0] _T_387 = {memRdata_flag_d,memRdata_flag_a,memRdata_flag_g,memRdata_flag_u,memRdata_flag_x,memRdata_flag_w,memRdata_flag_r,memRdata_flag_v}; // @[EmbeddedTLB.scala 292:44]
  wire  _T_398 = _T_387[1] | _T_387[3]; // @[EmbeddedTLB.scala 297:34]
  wire  _T_399 = ~_T_398; // @[EmbeddedTLB.scala 297:21]
  reg [1:0] level; // @[EmbeddedTLB.scala 248:22]
  wire  _T_400 = level == 2'h3; // @[EmbeddedTLB.scala 297:58]
  wire  _T_401 = level == 2'h2; // @[EmbeddedTLB.scala 297:73]
  wire  _T_402 = _T_400 | _T_401; // @[EmbeddedTLB.scala 297:65]
  wire  _T_403 = _T_399 & _T_402; // @[EmbeddedTLB.scala 297:49]
  wire  _T_404 = ~_T_387[0]; // @[EmbeddedTLB.scala 298:16]
  wire  _T_405 = ~_T_387[1]; // @[EmbeddedTLB.scala 298:32]
  wire  _T_406 = _T_405 & _T_387[2]; // @[EmbeddedTLB.scala 298:44]
  wire  _T_407 = _T_404 | _T_406; // @[EmbeddedTLB.scala 298:28]
  wire  _T_414 = _T_334 & _T_337; // @[EmbeddedTLB.scala 302:38]
  wire  _GEN_19 = _T_407 ? _T_414 : _T_338; // @[EmbeddedTLB.scala 298:60]
  wire  _T_451 = level != 2'h0; // @[EmbeddedTLB.scala 313:27]
  wire  _T_453 = ~_T_387[4]; // @[EmbeddedTLB.scala 314:74]
  wire  _T_454 = _T_314 & _T_453; // @[EmbeddedTLB.scala 314:71]
  wire  _T_455 = ~_T_454; // @[EmbeddedTLB.scala 314:41]
  wire  _T_456 = _T_387[0] & _T_455; // @[EmbeddedTLB.scala 314:38]
  wire  _T_458 = _T_319 & _T_387[4]; // @[EmbeddedTLB.scala 314:120]
  wire  _T_461 = _T_458 & _T_321; // @[EmbeddedTLB.scala 314:134]
  wire  _T_462 = ~_T_461; // @[EmbeddedTLB.scala 314:90]
  wire  _T_463 = _T_456 & _T_462; // @[EmbeddedTLB.scala 314:87]
  wire  _T_465 = io_pf_status_mxr & _T_387[3]; // @[EmbeddedTLB.scala 316:68]
  wire  _T_466 = _T_387[1] | _T_465; // @[EmbeddedTLB.scala 316:51]
  wire  _T_467 = _T_463 & _T_466; // @[EmbeddedTLB.scala 316:36]
  wire  _T_490 = ~_T_467; // @[EmbeddedTLB.scala 330:19]
  wire  _T_496 = _T_490 & _T_334; // @[EmbeddedTLB.scala 330:29]
  wire  _T_468 = _T_463 & _T_387[2]; // @[EmbeddedTLB.scala 317:37]
  wire  _T_497 = ~_T_468; // @[EmbeddedTLB.scala 330:50]
  wire  _T_499 = _T_497 & io_in_bits_cmd[0]; // @[EmbeddedTLB.scala 330:61]
  wire  _T_500 = _T_496 | _T_499; // @[EmbeddedTLB.scala 330:46]
  wire  _GEN_23 = _T_500 ? _T_414 : _T_338; // @[EmbeddedTLB.scala 330:80]
  wire  _GEN_29 = _T_451 ? _GEN_23 : _T_338; // @[EmbeddedTLB.scala 313:36]
  wire  _GEN_35 = _T_403 ? _GEN_19 : _GEN_29; // @[EmbeddedTLB.scala 297:82]
  wire  _GEN_54 = _T_397 ? _GEN_35 : _T_338; // @[EmbeddedTLB.scala 293:33]
  wire  _GEN_78 = _T_379 ? _GEN_54 : _T_338; // @[Conditional.scala 39:67]
  wire  _GEN_91 = _T_377 ? _T_338 : _GEN_78; // @[Conditional.scala 39:67]
  wire  loadPF = _T_370 ? _T_338 : _GEN_91; // @[Conditional.scala 40:58]
  wire  hitStore = hitCheck & hitFlag_w; // @[EmbeddedTLB.scala 229:27]
  wire  _T_339 = ~hitStore; // @[EmbeddedTLB.scala 242:17]
  wire  _T_341 = _T_339 & io_in_bits_cmd[0]; // @[EmbeddedTLB.scala 242:27]
  wire  _T_342 = _T_341 & hit; // @[EmbeddedTLB.scala 242:44]
  wire  _T_351 = _T_336 & ISAMO; // @[EmbeddedTLB.scala 242:88]
  wire  _T_352 = _T_342 | _T_351; // @[EmbeddedTLB.scala 242:52]
  wire  _T_416 = io_in_bits_cmd[0] | ISAMO; // @[EmbeddedTLB.scala 303:40]
  wire  _GEN_20 = _T_407 ? _T_416 : _T_352; // @[EmbeddedTLB.scala 298:60]
  wire  _GEN_24 = _T_500 ? _T_416 : _T_352; // @[EmbeddedTLB.scala 330:80]
  wire  _GEN_30 = _T_451 ? _GEN_24 : _T_352; // @[EmbeddedTLB.scala 313:36]
  wire  _GEN_36 = _T_403 ? _GEN_20 : _GEN_30; // @[EmbeddedTLB.scala 297:82]
  wire  _GEN_55 = _T_397 ? _GEN_36 : _T_352; // @[EmbeddedTLB.scala 293:33]
  wire  _GEN_79 = _T_379 ? _GEN_55 : _T_352; // @[Conditional.scala 39:67]
  wire  _GEN_92 = _T_377 ? _T_352 : _GEN_79; // @[Conditional.scala 39:67]
  wire  storePF = _T_370 ? _T_352 : _GEN_92; // @[Conditional.scala 40:58]
  wire  _T_297 = loadPF | storePF; // @[EmbeddedTLB.scala 221:93]
  wire  _T_298 = io_pf_loadPF | io_pf_storePF; // @[Bundle.scala 129:23]
  wire  _T_299 = _T_297 | _T_298; // @[EmbeddedTLB.scala 221:104]
  wire  _T_300 = ~_T_299; // @[EmbeddedTLB.scala 221:84]
  wire  hitWB = _T_294 & _T_300; // @[EmbeddedTLB.scala 221:81]
  wire [7:0] _T_303 = {io_in_bits_cmd[0],1'h1,6'h0}; // @[Cat.scala 29:58]
  wire [7:0] _T_310 = {hitFlag_d,hitFlag_a,hitFlag_g,hitFlag_u,hitFlag_x,hitFlag_w,hitFlag_r,hitFlag_v}; // @[EmbeddedTLB.scala 222:79]
  wire [7:0] hitRefillFlag = _T_303 | _T_310; // @[EmbeddedTLB.scala 222:69]
  wire [39:0] _T_313 = {10'h0,hitData_ppn,2'h0,hitRefillFlag}; // @[Cat.scala 29:58]
  reg [39:0] hitWBStore; // @[Reg.scala 15:16]
  reg  _T_327; // @[EmbeddedTLB.scala 236:26]
  reg  _T_328; // @[EmbeddedTLB.scala 237:27]
  reg [63:0] memRespStore; // @[EmbeddedTLB.scala 250:25]
  reg [17:0] missMaskStore; // @[EmbeddedTLB.scala 252:26]
  wire [19:0] memRdata_ppn = io_mem_resp_bits_rdata[29:10]; // @[EmbeddedTLB.scala 255:49]
  reg [31:0] raddr; // @[EmbeddedTLB.scala 256:18]
  wire  _T_365 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  reg  alreadyOutFire; // @[Reg.scala 27:20]
  wire  _GEN_2 = _T_365 | alreadyOutFire; // @[Reg.scala 28:19]
  wire [31:0] _T_376 = {satp_ppn,vpn_vpn2,3'h0}; // @[Cat.scala 29:58]
  wire  _T_378 = io_mem_req_ready & io_mem_req_valid; // @[Decoupled.scala 40:37]
  wire [8:0] _T_448 = _T_400 ? vpn_vpn1 : vpn_vpn0; // @[EmbeddedTLB.scala 311:50]
  wire [31:0] _T_450 = {memRdata_ppn,_T_448,3'h0}; // @[Cat.scala 29:58]
  wire  _T_469 = ~_T_387[6]; // @[EmbeddedTLB.scala 318:60]
  wire  _T_470 = ~_T_387[7]; // @[EmbeddedTLB.scala 318:76]
  wire  _T_472 = _T_470 & io_in_bits_cmd[0]; // @[EmbeddedTLB.scala 318:88]
  wire  _T_473 = _T_469 | _T_472; // @[EmbeddedTLB.scala 318:72]
  wire [63:0] _T_477 = {56'h0,io_in_bits_cmd[0],7'h40}; // @[Cat.scala 29:58]
  wire [7:0] _T_487 = {_T_387[7],_T_387[6],_T_387[5],_T_387[4],_T_387[3],_T_387[2],_T_387[1],_T_387[0]}; // @[EmbeddedTLB.scala 320:79]
  wire [7:0] _T_488 = _T_303 | _T_487; // @[EmbeddedTLB.scala 320:68]
  wire [63:0] _T_489 = io_mem_resp_bits_rdata | _T_477; // @[EmbeddedTLB.scala 321:50]
  wire  _GEN_25 = _T_500 ? 1'h0 : 1'h1; // @[EmbeddedTLB.scala 330:80]
  wire  _GEN_31 = _T_451 & _GEN_25; // @[EmbeddedTLB.scala 313:36]
  wire  _GEN_40 = _T_403 ? 1'h0 : _GEN_31; // @[EmbeddedTLB.scala 297:82]
  wire [1:0] _T_516 = level - 2'h1; // @[EmbeddedTLB.scala 342:24]
  wire  _GEN_59 = _T_397 & _GEN_40; // @[EmbeddedTLB.scala 293:33]
  wire  _T_517 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_519 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_523 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire  _GEN_83 = _T_379 & _GEN_59; // @[Conditional.scala 39:67]
  wire  _GEN_96 = _T_377 ? 1'h0 : _GEN_83; // @[Conditional.scala 39:67]
  wire  missMetaRefill = _T_370 ? 1'h0 : _GEN_96; // @[Conditional.scala 40:58]
  wire  cmd = state == 3'h3; // @[EmbeddedTLB.scala 365:23]
  wire  _T_527 = state == 3'h1; // @[EmbeddedTLB.scala 367:31]
  wire  _T_534 = state == 3'h0; // @[EmbeddedTLB.scala 371:82]
  wire  _T_535 = hitWB & _T_534; // @[EmbeddedTLB.scala 371:73]
  wire  _T_538 = missMetaRefill | _T_535; // @[EmbeddedTLB.scala 371:63]
  reg  _T_539; // @[EmbeddedTLB.scala 371:33]
  reg [3:0] _T_545; // @[EmbeddedTLB.scala 372:21]
  reg [3:0] _T_546; // @[EmbeddedTLB.scala 372:60]
  reg [26:0] _T_549; // @[EmbeddedTLB.scala 372:84]
  reg [15:0] _T_551; // @[EmbeddedTLB.scala 373:19]
  reg [17:0] _T_553; // @[EmbeddedTLB.scala 373:72]
  reg [7:0] _T_555; // @[EmbeddedTLB.scala 374:19]
  reg [19:0] _T_557; // @[EmbeddedTLB.scala 374:77]
  reg [31:0] _T_559; // @[EmbeddedTLB.scala 375:22]
  wire [59:0] _T_561 = {_T_555,_T_557,_T_559}; // @[Cat.scala 29:58]
  wire [60:0] _T_563 = {_T_549,_T_551,_T_553}; // @[Cat.scala 29:58]
  wire [31:0] _T_566 = {hitData_ppn,12'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_569 = {2'h3,hitMeta_mask,12'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_570 = _T_566 & _T_569; // @[BitUtils.scala 32:13]
  wire [31:0] _T_571 = ~_T_569; // @[BitUtils.scala 32:38]
  wire [31:0] _T_572 = io_in_bits_addr[31:0] & _T_571; // @[BitUtils.scala 32:36]
  wire [31:0] _T_573 = _T_570 | _T_572; // @[BitUtils.scala 32:25]
  wire [31:0] _T_588 = {memRespStore[29:10],12'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_591 = {2'h3,missMaskStore,12'h0}; // @[Cat.scala 29:58]
  wire [31:0] _T_592 = _T_588 & _T_591; // @[BitUtils.scala 32:13]
  wire [31:0] _T_593 = ~_T_591; // @[BitUtils.scala 32:38]
  wire [31:0] _T_594 = io_in_bits_addr[31:0] & _T_593; // @[BitUtils.scala 32:36]
  wire [31:0] _T_595 = _T_592 | _T_594; // @[BitUtils.scala 32:25]
  wire  _T_597 = ~hitWB; // @[EmbeddedTLB.scala 380:45]
  wire  _T_598 = hit & _T_597; // @[EmbeddedTLB.scala 380:42]
  wire  _T_600 = _T_298 | loadPF; // @[EmbeddedTLB.scala 380:68]
  wire  _T_601 = _T_600 | storePF; // @[EmbeddedTLB.scala 380:78]
  wire  _T_602 = ~_T_601; // @[EmbeddedTLB.scala 380:53]
  wire  _T_603 = state == 3'h4; // @[EmbeddedTLB.scala 380:97]
  wire  _T_604 = _T_598 ? _T_602 : _T_603; // @[EmbeddedTLB.scala 380:37]
  wire  _T_607 = io_out_ready & _T_534; // @[EmbeddedTLB.scala 382:31]
  wire  _T_608 = ~miss; // @[EmbeddedTLB.scala 382:56]
  wire  _T_609 = _T_607 & _T_608; // @[EmbeddedTLB.scala 382:53]
  wire  _T_611 = _T_609 & _T_597; // @[EmbeddedTLB.scala 382:62]
  wire  _T_612 = _T_611 & io_mdReady; // @[EmbeddedTLB.scala 382:72]
  wire  _T_614 = ~_T_298; // @[EmbeddedTLB.scala 382:90]
  wire  _T_615 = ~loadPF; // @[EmbeddedTLB.scala 382:107]
  wire  _T_616 = _T_614 & _T_615; // @[EmbeddedTLB.scala 382:104]
  wire  _T_617 = ~storePF; // @[EmbeddedTLB.scala 382:118]
  wire  _T_618 = _T_616 & _T_617; // @[EmbeddedTLB.scala 382:115]
  assign io_in_ready = _T_612 & _T_618; // @[EmbeddedTLB.scala 382:15]
  assign io_out_valid = io_in_valid & _T_604; // @[EmbeddedTLB.scala 380:16]
  assign io_out_bits_addr = hit ? _T_573 : _T_595; // @[EmbeddedTLB.scala 378:15 EmbeddedTLB.scala 379:20]
  assign io_out_bits_size = io_in_bits_size; // @[EmbeddedTLB.scala 378:15]
  assign io_out_bits_cmd = io_in_bits_cmd; // @[EmbeddedTLB.scala 378:15]
  assign io_out_bits_wmask = io_in_bits_wmask; // @[EmbeddedTLB.scala 378:15]
  assign io_out_bits_wdata = io_in_bits_wdata; // @[EmbeddedTLB.scala 378:15]
  assign io_mdWrite_wen = _T_539; // @[TLB.scala 214:14]
  assign io_mdWrite_windex = _T_545; // @[TLB.scala 215:17]
  assign io_mdWrite_waymask = _T_546; // @[TLB.scala 216:18]
  assign io_mdWrite_wdata = {_T_563,_T_561}; // @[TLB.scala 217:16]
  assign io_mem_req_valid = _T_527 | cmd; // @[EmbeddedTLB.scala 367:20]
  assign io_mem_req_bits_addr = hitWB ? hitData_pteaddr : raddr; // @[SimpleBus.scala 64:15]
  assign io_mem_req_bits_cmd = {{3'd0}, cmd}; // @[SimpleBus.scala 65:14]
  assign io_mem_req_bits_wdata = hitWB ? {{24'd0}, hitWBStore} : memRespStore; // @[SimpleBus.scala 67:16]
  assign io_mem_resp_ready = 1'h1; // @[EmbeddedTLB.scala 368:21]
  assign io_pf_loadPF = _T_327; // @[EmbeddedTLB.scala 199:13 EmbeddedTLB.scala 236:16]
  assign io_pf_storePF = _T_328; // @[EmbeddedTLB.scala 200:14 EmbeddedTLB.scala 237:17]
  assign io_pf_addr = io_in_bits_addr; // @[EmbeddedTLB.scala 201:11]
  assign io_isFinish = _T_365 | _T_298; // @[EmbeddedTLB.scala 385:15]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _T_227 = _RAND_0[63:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[2:0];
  _RAND_2 = {1{`RANDOM}};
  level = _RAND_2[1:0];
  _RAND_3 = {2{`RANDOM}};
  hitWBStore = _RAND_3[39:0];
  _RAND_4 = {1{`RANDOM}};
  _T_327 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_328 = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  memRespStore = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  missMaskStore = _RAND_7[17:0];
  _RAND_8 = {1{`RANDOM}};
  raddr = _RAND_8[31:0];
  _RAND_9 = {1{`RANDOM}};
  alreadyOutFire = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _T_539 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_545 = _RAND_11[3:0];
  _RAND_12 = {1{`RANDOM}};
  _T_546 = _RAND_12[3:0];
  _RAND_13 = {1{`RANDOM}};
  _T_549 = _RAND_13[26:0];
  _RAND_14 = {1{`RANDOM}};
  _T_551 = _RAND_14[15:0];
  _RAND_15 = {1{`RANDOM}};
  _T_553 = _RAND_15[17:0];
  _RAND_16 = {1{`RANDOM}};
  _T_555 = _RAND_16[7:0];
  _RAND_17 = {1{`RANDOM}};
  _T_557 = _RAND_17[19:0];
  _RAND_18 = {1{`RANDOM}};
  _T_559 = _RAND_18[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_227 <= 64'h1234567887654321;
    end else if (_T_235) begin
      _T_227 <= 64'h1;
    end else begin
      _T_227 <= _T_237;
    end
    if (reset) begin
      state <= 3'h0;
    end else if (_T_370) begin
      if (hitWB) begin
        state <= 3'h3;
      end else if (miss) begin
        state <= 3'h1;
      end
    end else if (_T_377) begin
      if (_T_378) begin
        state <= 3'h2;
      end
    end else if (_T_379) begin
      if (_T_397) begin
        if (_T_403) begin
          if (_T_407) begin
            state <= 3'h5;
          end else begin
            state <= 3'h1;
          end
        end else if (_T_451) begin
          if (_T_500) begin
            state <= 3'h5;
          end else if (_T_473) begin
            state <= 3'h3;
          end else begin
            state <= 3'h4;
          end
        end
      end
    end else if (_T_517) begin
      if (_T_378) begin
        state <= 3'h4;
      end
    end else if (_T_519) begin
      if (_GEN_2) begin
        state <= 3'h0;
      end
    end else if (_T_523) begin
      state <= 3'h0;
    end
    if (reset) begin
      level <= 2'h3;
    end else if (_T_370) begin
      if (!(hitWB)) begin
        if (miss) begin
          level <= 2'h3;
        end
      end
    end else if (!(_T_377)) begin
      if (_T_379) begin
        if (_T_397) begin
          level <= _T_516;
        end
      end
    end
    if (hitWB) begin
      hitWBStore <= _T_313;
    end
    if (reset) begin
      _T_327 <= 1'h0;
    end else if (_T_370) begin
      _T_327 <= _T_338;
    end else if (_T_377) begin
      _T_327 <= _T_338;
    end else if (_T_379) begin
      if (_T_397) begin
        if (_T_403) begin
          if (_T_407) begin
            _T_327 <= _T_414;
          end else begin
            _T_327 <= _T_338;
          end
        end else if (_T_451) begin
          if (_T_500) begin
            _T_327 <= _T_414;
          end else begin
            _T_327 <= _T_338;
          end
        end else begin
          _T_327 <= _T_338;
        end
      end else begin
        _T_327 <= _T_338;
      end
    end else begin
      _T_327 <= _T_338;
    end
    if (reset) begin
      _T_328 <= 1'h0;
    end else if (_T_370) begin
      _T_328 <= _T_352;
    end else if (_T_377) begin
      _T_328 <= _T_352;
    end else if (_T_379) begin
      if (_T_397) begin
        if (_T_403) begin
          if (_T_407) begin
            _T_328 <= _T_416;
          end else begin
            _T_328 <= _T_352;
          end
        end else if (_T_451) begin
          if (_T_500) begin
            _T_328 <= _T_416;
          end else begin
            _T_328 <= _T_352;
          end
        end else begin
          _T_328 <= _T_352;
        end
      end else begin
        _T_328 <= _T_352;
      end
    end else begin
      _T_328 <= _T_352;
    end
    if (!(_T_370)) begin
      if (!(_T_377)) begin
        if (_T_379) begin
          if (_T_397) begin
            if (!(_T_403)) begin
              if (_T_451) begin
                memRespStore <= _T_489;
              end
            end
          end
        end
      end
    end
    if (!(_T_370)) begin
      if (!(_T_377)) begin
        if (_T_379) begin
          if (_T_397) begin
            if (!(_T_403)) begin
              if (_T_451) begin
                if (_T_370) begin
                  missMaskStore <= 18'h3ffff;
                end else if (_T_377) begin
                  missMaskStore <= 18'h3ffff;
                end else if (_T_379) begin
                  if (_T_397) begin
                    if (_T_403) begin
                      missMaskStore <= 18'h3ffff;
                    end else if (_T_451) begin
                      if (_T_400) begin
                        missMaskStore <= 18'h0;
                      end else if (_T_401) begin
                        missMaskStore <= 18'h3fe00;
                      end else begin
                        missMaskStore <= 18'h3ffff;
                      end
                    end else begin
                      missMaskStore <= 18'h3ffff;
                    end
                  end else begin
                    missMaskStore <= 18'h3ffff;
                  end
                end else begin
                  missMaskStore <= 18'h3ffff;
                end
              end
            end
          end
        end
      end
    end
    if (_T_370) begin
      if (!(hitWB)) begin
        if (miss) begin
          raddr <= _T_376;
        end
      end
    end else if (!(_T_377)) begin
      if (_T_379) begin
        if (_T_397) begin
          if (_T_403) begin
            if (!(_T_407)) begin
              raddr <= _T_450;
            end
          end
        end
      end
    end
    if (reset) begin
      alreadyOutFire <= 1'h0;
    end else if (_T_370) begin
      if (hitWB) begin
        alreadyOutFire <= 1'h0;
      end else if (miss) begin
        alreadyOutFire <= 1'h0;
      end else begin
        alreadyOutFire <= _GEN_2;
      end
    end else if (_T_377) begin
      alreadyOutFire <= _GEN_2;
    end else if (_T_379) begin
      alreadyOutFire <= _GEN_2;
    end else if (_T_517) begin
      alreadyOutFire <= _GEN_2;
    end else if (_T_519) begin
      if (_GEN_2) begin
        alreadyOutFire <= 1'h0;
      end else begin
        alreadyOutFire <= _GEN_2;
      end
    end else begin
      alreadyOutFire <= _GEN_2;
    end
    if (reset) begin
      _T_539 <= 1'h0;
    end else begin
      _T_539 <= _T_538;
    end
    _T_545 <= io_in_bits_addr[15:12];
    if (hit) begin
      _T_546 <= hitVec;
    end else begin
      _T_546 <= victimWaymask;
    end
    _T_549 <= {_T_57,vpn_vpn0};
    if (hitWB) begin
      _T_551 <= hitMeta_asid;
    end else begin
      _T_551 <= satp_asid;
    end
    if (hitWB) begin
      _T_553 <= hitMeta_mask;
    end else if (_T_370) begin
      _T_553 <= 18'h3ffff;
    end else if (_T_377) begin
      _T_553 <= 18'h3ffff;
    end else if (_T_379) begin
      if (_T_397) begin
        if (_T_403) begin
          _T_553 <= 18'h3ffff;
        end else if (_T_451) begin
          if (_T_400) begin
            _T_553 <= 18'h0;
          end else if (_T_401) begin
            _T_553 <= 18'h3fe00;
          end else begin
            _T_553 <= 18'h3ffff;
          end
        end else begin
          _T_553 <= 18'h3ffff;
        end
      end else begin
        _T_553 <= 18'h3ffff;
      end
    end else begin
      _T_553 <= 18'h3ffff;
    end
    if (hitWB) begin
      _T_555 <= hitRefillFlag;
    end else if (_T_370) begin
      _T_555 <= 8'h0;
    end else if (_T_377) begin
      _T_555 <= 8'h0;
    end else if (_T_379) begin
      if (_T_397) begin
        if (_T_403) begin
          _T_555 <= 8'h0;
        end else if (_T_451) begin
          _T_555 <= _T_488;
        end else begin
          _T_555 <= 8'h0;
        end
      end else begin
        _T_555 <= 8'h0;
      end
    end else begin
      _T_555 <= 8'h0;
    end
    if (hitWB) begin
      _T_557 <= hitData_ppn;
    end else begin
      _T_557 <= memRdata_ppn;
    end
    if (hitWB) begin
      _T_559 <= hitData_pteaddr;
    end else begin
      _T_559 <= raddr;
    end
  end
endmodule
module EmbeddedTLBEmpty_1(
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [2:0]  io_in_bits_size,
  input  [3:0]  io_in_bits_cmd,
  input  [7:0]  io_in_bits_wmask,
  input  [63:0] io_in_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [2:0]  io_out_bits_size,
  output [3:0]  io_out_bits_cmd,
  output [7:0]  io_out_bits_wmask,
  output [63:0] io_out_bits_wdata
);
  assign io_in_ready = io_out_ready; // @[EmbeddedTLB.scala 403:10]
  assign io_out_valid = io_in_valid; // @[EmbeddedTLB.scala 403:10]
  assign io_out_bits_addr = io_in_bits_addr; // @[EmbeddedTLB.scala 403:10]
  assign io_out_bits_size = io_in_bits_size; // @[EmbeddedTLB.scala 403:10]
  assign io_out_bits_cmd = io_in_bits_cmd; // @[EmbeddedTLB.scala 403:10]
  assign io_out_bits_wmask = io_in_bits_wmask; // @[EmbeddedTLB.scala 403:10]
  assign io_out_bits_wdata = io_in_bits_wdata; // @[EmbeddedTLB.scala 403:10]
endmodule
module EmbeddedTLBMD_1(
  input          clock,
  input          reset,
  output [120:0] io_tlbmd_0,
  output [120:0] io_tlbmd_1,
  output [120:0] io_tlbmd_2,
  output [120:0] io_tlbmd_3,
  input          io_write_wen,
  input  [3:0]   io_write_windex,
  input  [3:0]   io_write_waymask,
  input  [120:0] io_write_wdata,
  input  [3:0]   io_rindex,
  output         io_ready
);
`ifdef RANDOMIZE_MEM_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [120:0] tlbmd_0 [0:15]; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_0__T_data; // @[EmbeddedTLB.scala 38:18]
  wire [3:0] tlbmd_0__T_addr; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_0__T_9_data; // @[EmbeddedTLB.scala 38:18]
  wire [3:0] tlbmd_0__T_9_addr; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_0__T_9_mask; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_0__T_9_en; // @[EmbeddedTLB.scala 38:18]
  reg [120:0] tlbmd_1 [0:15]; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_1__T_data; // @[EmbeddedTLB.scala 38:18]
  wire [3:0] tlbmd_1__T_addr; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_1__T_9_data; // @[EmbeddedTLB.scala 38:18]
  wire [3:0] tlbmd_1__T_9_addr; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_1__T_9_mask; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_1__T_9_en; // @[EmbeddedTLB.scala 38:18]
  reg [120:0] tlbmd_2 [0:15]; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_2__T_data; // @[EmbeddedTLB.scala 38:18]
  wire [3:0] tlbmd_2__T_addr; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_2__T_9_data; // @[EmbeddedTLB.scala 38:18]
  wire [3:0] tlbmd_2__T_9_addr; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_2__T_9_mask; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_2__T_9_en; // @[EmbeddedTLB.scala 38:18]
  reg [120:0] tlbmd_3 [0:15]; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_3__T_data; // @[EmbeddedTLB.scala 38:18]
  wire [3:0] tlbmd_3__T_addr; // @[EmbeddedTLB.scala 38:18]
  wire [120:0] tlbmd_3__T_9_data; // @[EmbeddedTLB.scala 38:18]
  wire [3:0] tlbmd_3__T_9_addr; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_3__T_9_mask; // @[EmbeddedTLB.scala 38:18]
  wire  tlbmd_3__T_9_en; // @[EmbeddedTLB.scala 38:18]
  reg  resetState; // @[EmbeddedTLB.scala 42:27]
  reg [3:0] resetSet; // @[Counter.scala 29:33]
  wire  _T_1 = resetSet == 4'hf; // @[Counter.scala 38:24]
  wire [3:0] _T_3 = resetSet + 4'h1; // @[Counter.scala 39:22]
  wire  resetFinish = resetState & _T_1; // @[Counter.scala 67:17]
  wire  _GEN_2 = resetFinish ? 1'h0 : resetState; // @[EmbeddedTLB.scala 44:22]
  wire [3:0] waymask = resetState ? 4'hf : io_write_waymask; // @[EmbeddedTLB.scala 53:20]
  assign tlbmd_0__T_addr = io_rindex;
  assign tlbmd_0__T_data = tlbmd_0[tlbmd_0__T_addr]; // @[EmbeddedTLB.scala 38:18]
  assign tlbmd_0__T_9_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_0__T_9_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_0__T_9_mask = waymask[0];
  assign tlbmd_0__T_9_en = resetState | io_write_wen;
  assign tlbmd_1__T_addr = io_rindex;
  assign tlbmd_1__T_data = tlbmd_1[tlbmd_1__T_addr]; // @[EmbeddedTLB.scala 38:18]
  assign tlbmd_1__T_9_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_1__T_9_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_1__T_9_mask = waymask[1];
  assign tlbmd_1__T_9_en = resetState | io_write_wen;
  assign tlbmd_2__T_addr = io_rindex;
  assign tlbmd_2__T_data = tlbmd_2[tlbmd_2__T_addr]; // @[EmbeddedTLB.scala 38:18]
  assign tlbmd_2__T_9_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_2__T_9_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_2__T_9_mask = waymask[2];
  assign tlbmd_2__T_9_en = resetState | io_write_wen;
  assign tlbmd_3__T_addr = io_rindex;
  assign tlbmd_3__T_data = tlbmd_3[tlbmd_3__T_addr]; // @[EmbeddedTLB.scala 38:18]
  assign tlbmd_3__T_9_data = resetState ? 121'h0 : io_write_wdata;
  assign tlbmd_3__T_9_addr = resetState ? resetSet : io_write_windex;
  assign tlbmd_3__T_9_mask = waymask[3];
  assign tlbmd_3__T_9_en = resetState | io_write_wen;
  assign io_tlbmd_0 = tlbmd_0__T_data; // @[EmbeddedTLB.scala 39:12]
  assign io_tlbmd_1 = tlbmd_1__T_data; // @[EmbeddedTLB.scala 39:12]
  assign io_tlbmd_2 = tlbmd_2__T_data; // @[EmbeddedTLB.scala 39:12]
  assign io_tlbmd_3 = tlbmd_3__T_data; // @[EmbeddedTLB.scala 39:12]
  assign io_ready = ~resetState; // @[EmbeddedTLB.scala 59:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {4{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_0[initvar] = _RAND_0[120:0];
  _RAND_1 = {4{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_1[initvar] = _RAND_1[120:0];
  _RAND_2 = {4{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_2[initvar] = _RAND_2[120:0];
  _RAND_3 = {4{`RANDOM}};
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    tlbmd_3[initvar] = _RAND_3[120:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  resetState = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  resetSet = _RAND_5[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(tlbmd_0__T_9_en & tlbmd_0__T_9_mask) begin
      tlbmd_0[tlbmd_0__T_9_addr] <= tlbmd_0__T_9_data; // @[EmbeddedTLB.scala 38:18]
    end
    if(tlbmd_1__T_9_en & tlbmd_1__T_9_mask) begin
      tlbmd_1[tlbmd_1__T_9_addr] <= tlbmd_1__T_9_data; // @[EmbeddedTLB.scala 38:18]
    end
    if(tlbmd_2__T_9_en & tlbmd_2__T_9_mask) begin
      tlbmd_2[tlbmd_2__T_9_addr] <= tlbmd_2__T_9_data; // @[EmbeddedTLB.scala 38:18]
    end
    if(tlbmd_3__T_9_en & tlbmd_3__T_9_mask) begin
      tlbmd_3[tlbmd_3__T_9_addr] <= tlbmd_3__T_9_data; // @[EmbeddedTLB.scala 38:18]
    end
    resetState <= reset | _GEN_2;
    if (reset) begin
      resetSet <= 4'h0;
    end else if (resetState) begin
      resetSet <= _T_3;
    end
  end
endmodule
module EmbeddedTLB_1(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [38:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [2:0]  io_out_req_bits_size,
  output [3:0]  io_out_req_bits_cmd,
  output [7:0]  io_out_req_bits_wmask,
  output [63:0] io_out_req_bits_wdata,
  input         io_out_resp_valid,
  input  [63:0] io_out_resp_bits_rdata,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [31:0] io_mem_req_bits_addr,
  output [3:0]  io_mem_req_bits_cmd,
  output [63:0] io_mem_req_bits_wdata,
  input         io_mem_resp_valid,
  input  [63:0] io_mem_resp_bits_rdata,
  input  [1:0]  io_csrMMU_priviledgeMode,
  input         io_csrMMU_status_sum,
  input         io_csrMMU_status_mxr,
  output        io_csrMMU_loadPF,
  output        io_csrMMU_storePF,
  output [38:0] io_csrMMU_addr,
  output        _T_38_0,
  input  [63:0] CSRSATP,
  input         amoReq,
  output        vmEnable_0,
  output        _T_37_0,
  input         MOUFlushTLB
);
`ifdef RANDOMIZE_REG_INIT
  reg [127:0] _RAND_0;
  reg [127:0] _RAND_1;
  reg [127:0] _RAND_2;
  reg [127:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [63:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  tlbExec_clock; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_reset; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_in_ready; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_in_valid; // @[EmbeddedTLB.scala 80:23]
  wire [38:0] tlbExec_io_in_bits_addr; // @[EmbeddedTLB.scala 80:23]
  wire [2:0] tlbExec_io_in_bits_size; // @[EmbeddedTLB.scala 80:23]
  wire [3:0] tlbExec_io_in_bits_cmd; // @[EmbeddedTLB.scala 80:23]
  wire [7:0] tlbExec_io_in_bits_wmask; // @[EmbeddedTLB.scala 80:23]
  wire [63:0] tlbExec_io_in_bits_wdata; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_out_ready; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_out_valid; // @[EmbeddedTLB.scala 80:23]
  wire [31:0] tlbExec_io_out_bits_addr; // @[EmbeddedTLB.scala 80:23]
  wire [2:0] tlbExec_io_out_bits_size; // @[EmbeddedTLB.scala 80:23]
  wire [3:0] tlbExec_io_out_bits_cmd; // @[EmbeddedTLB.scala 80:23]
  wire [7:0] tlbExec_io_out_bits_wmask; // @[EmbeddedTLB.scala 80:23]
  wire [63:0] tlbExec_io_out_bits_wdata; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_md_0; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_md_1; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_md_2; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_md_3; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mdWrite_wen; // @[EmbeddedTLB.scala 80:23]
  wire [3:0] tlbExec_io_mdWrite_windex; // @[EmbeddedTLB.scala 80:23]
  wire [3:0] tlbExec_io_mdWrite_waymask; // @[EmbeddedTLB.scala 80:23]
  wire [120:0] tlbExec_io_mdWrite_wdata; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mdReady; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mem_req_ready; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mem_req_valid; // @[EmbeddedTLB.scala 80:23]
  wire [31:0] tlbExec_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 80:23]
  wire [3:0] tlbExec_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 80:23]
  wire [63:0] tlbExec_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mem_resp_ready; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_mem_resp_valid; // @[EmbeddedTLB.scala 80:23]
  wire [63:0] tlbExec_io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 80:23]
  wire [63:0] tlbExec_io_satp; // @[EmbeddedTLB.scala 80:23]
  wire [1:0] tlbExec_io_pf_priviledgeMode; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_pf_status_sum; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_pf_status_mxr; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_pf_loadPF; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_pf_storePF; // @[EmbeddedTLB.scala 80:23]
  wire [38:0] tlbExec_io_pf_addr; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_io_isFinish; // @[EmbeddedTLB.scala 80:23]
  wire  tlbExec_ISAMO; // @[EmbeddedTLB.scala 80:23]
  wire  tlbEmpty_io_in_ready; // @[EmbeddedTLB.scala 81:24]
  wire  tlbEmpty_io_in_valid; // @[EmbeddedTLB.scala 81:24]
  wire [31:0] tlbEmpty_io_in_bits_addr; // @[EmbeddedTLB.scala 81:24]
  wire [2:0] tlbEmpty_io_in_bits_size; // @[EmbeddedTLB.scala 81:24]
  wire [3:0] tlbEmpty_io_in_bits_cmd; // @[EmbeddedTLB.scala 81:24]
  wire [7:0] tlbEmpty_io_in_bits_wmask; // @[EmbeddedTLB.scala 81:24]
  wire [63:0] tlbEmpty_io_in_bits_wdata; // @[EmbeddedTLB.scala 81:24]
  wire  tlbEmpty_io_out_ready; // @[EmbeddedTLB.scala 81:24]
  wire  tlbEmpty_io_out_valid; // @[EmbeddedTLB.scala 81:24]
  wire [31:0] tlbEmpty_io_out_bits_addr; // @[EmbeddedTLB.scala 81:24]
  wire [2:0] tlbEmpty_io_out_bits_size; // @[EmbeddedTLB.scala 81:24]
  wire [3:0] tlbEmpty_io_out_bits_cmd; // @[EmbeddedTLB.scala 81:24]
  wire [7:0] tlbEmpty_io_out_bits_wmask; // @[EmbeddedTLB.scala 81:24]
  wire [63:0] tlbEmpty_io_out_bits_wdata; // @[EmbeddedTLB.scala 81:24]
  wire  mdTLB_clock; // @[EmbeddedTLB.scala 82:21]
  wire  mdTLB_reset; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_tlbmd_0; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_tlbmd_1; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_tlbmd_2; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_tlbmd_3; // @[EmbeddedTLB.scala 82:21]
  wire  mdTLB_io_write_wen; // @[EmbeddedTLB.scala 82:21]
  wire [3:0] mdTLB_io_write_windex; // @[EmbeddedTLB.scala 82:21]
  wire [3:0] mdTLB_io_write_waymask; // @[EmbeddedTLB.scala 82:21]
  wire [120:0] mdTLB_io_write_wdata; // @[EmbeddedTLB.scala 82:21]
  wire [3:0] mdTLB_io_rindex; // @[EmbeddedTLB.scala 82:21]
  wire  mdTLB_io_ready; // @[EmbeddedTLB.scala 82:21]
  reg [120:0] _T__0; // @[Reg.scala 15:16]
  reg [120:0] _T__1; // @[Reg.scala 15:16]
  reg [120:0] _T__2; // @[Reg.scala 15:16]
  reg [120:0] _T__3; // @[Reg.scala 15:16]
  wire  mdUpdate = io_in_req_valid & tlbExec_io_in_ready; // @[EmbeddedTLB.scala 114:26]
  wire  _T_14 = CSRSATP[63:60] == 4'h8; // @[EmbeddedTLB.scala 102:49]
  wire  _T_15 = io_csrMMU_priviledgeMode < 2'h3; // @[EmbeddedTLB.scala 102:86]
  wire  vmEnable = _T_14 & _T_15; // @[EmbeddedTLB.scala 102:57]
  reg  _T_16; // @[EmbeddedTLB.scala 105:24]
  wire  _GEN_4 = tlbExec_io_isFinish ? 1'h0 : _T_16; // @[EmbeddedTLB.scala 106:25]
  wire  _T_18 = mdUpdate & vmEnable; // @[EmbeddedTLB.scala 107:37]
  wire  _GEN_5 = _T_18 | _GEN_4; // @[EmbeddedTLB.scala 107:50]
  reg [38:0] _T_20_addr; // @[Reg.scala 15:16]
  reg [2:0] _T_20_size; // @[Reg.scala 15:16]
  reg [3:0] _T_20_cmd; // @[Reg.scala 15:16]
  reg [7:0] _T_20_wmask; // @[Reg.scala 15:16]
  reg [63:0] _T_20_wdata; // @[Reg.scala 15:16]
  wire  _T_22 = tlbEmpty_io_out_ready & tlbEmpty_io_out_valid; // @[Decoupled.scala 40:37]
  reg  _T_23; // @[Pipeline.scala 24:24]
  wire  _GEN_12 = _T_22 ? 1'h0 : _T_23; // @[Pipeline.scala 25:25]
  wire  _T_24 = tlbExec_io_out_valid & tlbEmpty_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_13 = _T_24 | _GEN_12; // @[Pipeline.scala 26:38]
  reg [31:0] _T_26_addr; // @[Reg.scala 15:16]
  reg [2:0] _T_26_size; // @[Reg.scala 15:16]
  reg [3:0] _T_26_cmd; // @[Reg.scala 15:16]
  reg [7:0] _T_26_wmask; // @[Reg.scala 15:16]
  reg [63:0] _T_26_wdata; // @[Reg.scala 15:16]
  wire  _T_27 = ~vmEnable; // @[EmbeddedTLB.scala 123:8]
  wire  _T_29 = ~tlbExec_io_out_ready; // @[EmbeddedTLB.scala 142:84]
  wire  _T_30 = tlbExec_io_out_valid & _T_29; // @[EmbeddedTLB.scala 142:81]
  reg  _T_31; // @[Reg.scala 27:20]
  wire  _GEN_29 = _T_30 | _T_31; // @[Reg.scala 28:19]
  wire  _T_32 = tlbExec_io_out_ready & tlbExec_io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_33 = _T_31 & _T_32; // @[EmbeddedTLB.scala 143:27]
  wire  _T_34 = ~_T_31; // @[EmbeddedTLB.scala 144:46]
  wire  _T_35 = tlbExec_io_out_valid & _T_34; // @[EmbeddedTLB.scala 144:43]
  wire  _T_36 = tlbExec_io_pf_loadPF | tlbExec_io_pf_storePF; // @[Bundle.scala 129:23]
  wire  _T_37 = _T_35 | _T_36; // @[EmbeddedTLB.scala 144:65]
  wire  _T_38 = io_csrMMU_loadPF | io_csrMMU_storePF; // @[Bundle.scala 129:23]
  EmbeddedTLBExec_1 tlbExec ( // @[EmbeddedTLB.scala 80:23]
    .clock(tlbExec_clock),
    .reset(tlbExec_reset),
    .io_in_ready(tlbExec_io_in_ready),
    .io_in_valid(tlbExec_io_in_valid),
    .io_in_bits_addr(tlbExec_io_in_bits_addr),
    .io_in_bits_size(tlbExec_io_in_bits_size),
    .io_in_bits_cmd(tlbExec_io_in_bits_cmd),
    .io_in_bits_wmask(tlbExec_io_in_bits_wmask),
    .io_in_bits_wdata(tlbExec_io_in_bits_wdata),
    .io_out_ready(tlbExec_io_out_ready),
    .io_out_valid(tlbExec_io_out_valid),
    .io_out_bits_addr(tlbExec_io_out_bits_addr),
    .io_out_bits_size(tlbExec_io_out_bits_size),
    .io_out_bits_cmd(tlbExec_io_out_bits_cmd),
    .io_out_bits_wmask(tlbExec_io_out_bits_wmask),
    .io_out_bits_wdata(tlbExec_io_out_bits_wdata),
    .io_md_0(tlbExec_io_md_0),
    .io_md_1(tlbExec_io_md_1),
    .io_md_2(tlbExec_io_md_2),
    .io_md_3(tlbExec_io_md_3),
    .io_mdWrite_wen(tlbExec_io_mdWrite_wen),
    .io_mdWrite_windex(tlbExec_io_mdWrite_windex),
    .io_mdWrite_waymask(tlbExec_io_mdWrite_waymask),
    .io_mdWrite_wdata(tlbExec_io_mdWrite_wdata),
    .io_mdReady(tlbExec_io_mdReady),
    .io_mem_req_ready(tlbExec_io_mem_req_ready),
    .io_mem_req_valid(tlbExec_io_mem_req_valid),
    .io_mem_req_bits_addr(tlbExec_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(tlbExec_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(tlbExec_io_mem_req_bits_wdata),
    .io_mem_resp_ready(tlbExec_io_mem_resp_ready),
    .io_mem_resp_valid(tlbExec_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(tlbExec_io_mem_resp_bits_rdata),
    .io_satp(tlbExec_io_satp),
    .io_pf_priviledgeMode(tlbExec_io_pf_priviledgeMode),
    .io_pf_status_sum(tlbExec_io_pf_status_sum),
    .io_pf_status_mxr(tlbExec_io_pf_status_mxr),
    .io_pf_loadPF(tlbExec_io_pf_loadPF),
    .io_pf_storePF(tlbExec_io_pf_storePF),
    .io_pf_addr(tlbExec_io_pf_addr),
    .io_isFinish(tlbExec_io_isFinish),
    .ISAMO(tlbExec_ISAMO)
  );
  EmbeddedTLBEmpty_1 tlbEmpty ( // @[EmbeddedTLB.scala 81:24]
    .io_in_ready(tlbEmpty_io_in_ready),
    .io_in_valid(tlbEmpty_io_in_valid),
    .io_in_bits_addr(tlbEmpty_io_in_bits_addr),
    .io_in_bits_size(tlbEmpty_io_in_bits_size),
    .io_in_bits_cmd(tlbEmpty_io_in_bits_cmd),
    .io_in_bits_wmask(tlbEmpty_io_in_bits_wmask),
    .io_in_bits_wdata(tlbEmpty_io_in_bits_wdata),
    .io_out_ready(tlbEmpty_io_out_ready),
    .io_out_valid(tlbEmpty_io_out_valid),
    .io_out_bits_addr(tlbEmpty_io_out_bits_addr),
    .io_out_bits_size(tlbEmpty_io_out_bits_size),
    .io_out_bits_cmd(tlbEmpty_io_out_bits_cmd),
    .io_out_bits_wmask(tlbEmpty_io_out_bits_wmask),
    .io_out_bits_wdata(tlbEmpty_io_out_bits_wdata)
  );
  EmbeddedTLBMD_1 mdTLB ( // @[EmbeddedTLB.scala 82:21]
    .clock(mdTLB_clock),
    .reset(mdTLB_reset),
    .io_tlbmd_0(mdTLB_io_tlbmd_0),
    .io_tlbmd_1(mdTLB_io_tlbmd_1),
    .io_tlbmd_2(mdTLB_io_tlbmd_2),
    .io_tlbmd_3(mdTLB_io_tlbmd_3),
    .io_write_wen(mdTLB_io_write_wen),
    .io_write_windex(mdTLB_io_write_windex),
    .io_write_waymask(mdTLB_io_write_waymask),
    .io_write_wdata(mdTLB_io_write_wdata),
    .io_rindex(mdTLB_io_rindex),
    .io_ready(mdTLB_io_ready)
  );
  assign io_in_req_ready = _T_27 ? io_out_req_ready : tlbExec_io_in_ready; // @[EmbeddedTLB.scala 110:16 EmbeddedTLB.scala 127:21]
  assign io_in_resp_valid = io_out_resp_valid; // @[EmbeddedTLB.scala 138:15]
  assign io_in_resp_bits_rdata = io_out_resp_bits_rdata; // @[EmbeddedTLB.scala 138:15]
  assign io_out_req_valid = _T_27 ? io_in_req_valid : tlbEmpty_io_out_valid; // @[EmbeddedTLB.scala 126:22 EmbeddedTLB.scala 135:41]
  assign io_out_req_bits_addr = _T_27 ? io_in_req_bits_addr[31:0] : tlbEmpty_io_out_bits_addr; // @[EmbeddedTLB.scala 128:26 EmbeddedTLB.scala 135:41]
  assign io_out_req_bits_size = _T_27 ? io_in_req_bits_size : tlbEmpty_io_out_bits_size; // @[EmbeddedTLB.scala 129:26 EmbeddedTLB.scala 135:41]
  assign io_out_req_bits_cmd = _T_27 ? io_in_req_bits_cmd : tlbEmpty_io_out_bits_cmd; // @[EmbeddedTLB.scala 130:25 EmbeddedTLB.scala 135:41]
  assign io_out_req_bits_wmask = _T_27 ? io_in_req_bits_wmask : tlbEmpty_io_out_bits_wmask; // @[EmbeddedTLB.scala 131:27 EmbeddedTLB.scala 135:41]
  assign io_out_req_bits_wdata = _T_27 ? io_in_req_bits_wdata : tlbEmpty_io_out_bits_wdata; // @[EmbeddedTLB.scala 132:27 EmbeddedTLB.scala 135:41]
  assign io_mem_req_valid = tlbExec_io_mem_req_valid; // @[EmbeddedTLB.scala 87:18]
  assign io_mem_req_bits_addr = tlbExec_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 87:18]
  assign io_mem_req_bits_cmd = tlbExec_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 87:18]
  assign io_mem_req_bits_wdata = tlbExec_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 87:18]
  assign io_csrMMU_loadPF = tlbExec_io_pf_loadPF; // @[EmbeddedTLB.scala 88:17]
  assign io_csrMMU_storePF = tlbExec_io_pf_storePF; // @[EmbeddedTLB.scala 88:17]
  assign io_csrMMU_addr = tlbExec_io_pf_addr; // @[EmbeddedTLB.scala 88:17]
  assign _T_38_0 = _T_38;
  assign vmEnable_0 = vmEnable;
  assign _T_37_0 = _T_37;
  assign tlbExec_clock = clock;
  assign tlbExec_reset = reset;
  assign tlbExec_io_in_valid = _T_16; // @[EmbeddedTLB.scala 112:17]
  assign tlbExec_io_in_bits_addr = _T_20_addr; // @[EmbeddedTLB.scala 111:16]
  assign tlbExec_io_in_bits_size = _T_20_size; // @[EmbeddedTLB.scala 111:16]
  assign tlbExec_io_in_bits_cmd = _T_20_cmd; // @[EmbeddedTLB.scala 111:16]
  assign tlbExec_io_in_bits_wmask = _T_20_wmask; // @[EmbeddedTLB.scala 111:16]
  assign tlbExec_io_in_bits_wdata = _T_20_wdata; // @[EmbeddedTLB.scala 111:16]
  assign tlbExec_io_out_ready = _T_27 | tlbEmpty_io_in_ready; // @[Pipeline.scala 29:16 EmbeddedTLB.scala 124:26]
  assign tlbExec_io_md_0 = _T__0; // @[EmbeddedTLB.scala 89:17]
  assign tlbExec_io_md_1 = _T__1; // @[EmbeddedTLB.scala 89:17]
  assign tlbExec_io_md_2 = _T__2; // @[EmbeddedTLB.scala 89:17]
  assign tlbExec_io_md_3 = _T__3; // @[EmbeddedTLB.scala 89:17]
  assign tlbExec_io_mdReady = mdTLB_io_ready; // @[EmbeddedTLB.scala 90:22]
  assign tlbExec_io_mem_req_ready = io_mem_req_ready; // @[EmbeddedTLB.scala 87:18]
  assign tlbExec_io_mem_resp_valid = io_mem_resp_valid; // @[EmbeddedTLB.scala 87:18]
  assign tlbExec_io_mem_resp_bits_rdata = io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 87:18]
  assign tlbExec_io_satp = CSRSATP; // @[EmbeddedTLB.scala 86:19]
  assign tlbExec_io_pf_priviledgeMode = io_csrMMU_priviledgeMode; // @[EmbeddedTLB.scala 88:17]
  assign tlbExec_io_pf_status_sum = io_csrMMU_status_sum; // @[EmbeddedTLB.scala 88:17]
  assign tlbExec_io_pf_status_mxr = io_csrMMU_status_mxr; // @[EmbeddedTLB.scala 88:17]
  assign tlbExec_ISAMO = amoReq;
  assign tlbEmpty_io_in_valid = _T_23; // @[Pipeline.scala 31:17]
  assign tlbEmpty_io_in_bits_addr = _T_26_addr; // @[Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_size = _T_26_size; // @[Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_cmd = _T_26_cmd; // @[Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_wmask = _T_26_wmask; // @[Pipeline.scala 30:16]
  assign tlbEmpty_io_in_bits_wdata = _T_26_wdata; // @[Pipeline.scala 30:16]
  assign tlbEmpty_io_out_ready = _T_27 | io_out_req_ready; // @[EmbeddedTLB.scala 125:52 EmbeddedTLB.scala 135:41]
  assign mdTLB_clock = clock;
  assign mdTLB_reset = reset | MOUFlushTLB; // @[EmbeddedTLB.scala 99:15]
  assign mdTLB_io_write_wen = tlbExec_io_mdWrite_wen; // @[EmbeddedTLB.scala 92:18]
  assign mdTLB_io_write_windex = tlbExec_io_mdWrite_windex; // @[EmbeddedTLB.scala 92:18]
  assign mdTLB_io_write_waymask = tlbExec_io_mdWrite_waymask; // @[EmbeddedTLB.scala 92:18]
  assign mdTLB_io_write_wdata = tlbExec_io_mdWrite_wdata; // @[EmbeddedTLB.scala 92:18]
  assign mdTLB_io_rindex = io_in_req_bits_addr[15:12]; // @[EmbeddedTLB.scala 91:19]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {4{`RANDOM}};
  _T__0 = _RAND_0[120:0];
  _RAND_1 = {4{`RANDOM}};
  _T__1 = _RAND_1[120:0];
  _RAND_2 = {4{`RANDOM}};
  _T__2 = _RAND_2[120:0];
  _RAND_3 = {4{`RANDOM}};
  _T__3 = _RAND_3[120:0];
  _RAND_4 = {1{`RANDOM}};
  _T_16 = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  _T_20_addr = _RAND_5[38:0];
  _RAND_6 = {1{`RANDOM}};
  _T_20_size = _RAND_6[2:0];
  _RAND_7 = {1{`RANDOM}};
  _T_20_cmd = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  _T_20_wmask = _RAND_8[7:0];
  _RAND_9 = {2{`RANDOM}};
  _T_20_wdata = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  _T_23 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_26_addr = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  _T_26_size = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  _T_26_cmd = _RAND_13[3:0];
  _RAND_14 = {1{`RANDOM}};
  _T_26_wmask = _RAND_14[7:0];
  _RAND_15 = {2{`RANDOM}};
  _T_26_wdata = _RAND_15[63:0];
  _RAND_16 = {1{`RANDOM}};
  _T_31 = _RAND_16[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (mdUpdate) begin
      _T__0 <= mdTLB_io_tlbmd_0;
    end
    if (mdUpdate) begin
      _T__1 <= mdTLB_io_tlbmd_1;
    end
    if (mdUpdate) begin
      _T__2 <= mdTLB_io_tlbmd_2;
    end
    if (mdUpdate) begin
      _T__3 <= mdTLB_io_tlbmd_3;
    end
    if (reset) begin
      _T_16 <= 1'h0;
    end else begin
      _T_16 <= _GEN_5;
    end
    if (mdUpdate) begin
      _T_20_addr <= io_in_req_bits_addr;
    end
    if (mdUpdate) begin
      _T_20_size <= io_in_req_bits_size;
    end
    if (mdUpdate) begin
      _T_20_cmd <= io_in_req_bits_cmd;
    end
    if (mdUpdate) begin
      _T_20_wmask <= io_in_req_bits_wmask;
    end
    if (mdUpdate) begin
      _T_20_wdata <= io_in_req_bits_wdata;
    end
    if (reset) begin
      _T_23 <= 1'h0;
    end else begin
      _T_23 <= _GEN_13;
    end
    if (_T_24) begin
      _T_26_addr <= tlbExec_io_out_bits_addr;
    end
    if (_T_24) begin
      _T_26_size <= tlbExec_io_out_bits_size;
    end
    if (_T_24) begin
      _T_26_cmd <= tlbExec_io_out_bits_cmd;
    end
    if (_T_24) begin
      _T_26_wmask <= tlbExec_io_out_bits_wmask;
    end
    if (_T_24) begin
      _T_26_wdata <= tlbExec_io_out_bits_wdata;
    end
    if (reset) begin
      _T_31 <= 1'h0;
    end else if (_T_33) begin
      _T_31 <= 1'h0;
    end else begin
      _T_31 <= _GEN_29;
    end
  end
endmodule
module CacheStage1_1(
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [2:0]  io_in_bits_size,
  input  [3:0]  io_in_bits_cmd,
  input  [7:0]  io_in_bits_wmask,
  input  [63:0] io_in_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [2:0]  io_out_bits_req_size,
  output [3:0]  io_out_bits_req_cmd,
  output [7:0]  io_out_bits_req_wmask,
  output [63:0] io_out_bits_req_wdata,
  input         io_metaReadBus_req_ready,
  output        io_metaReadBus_req_valid,
  output [6:0]  io_metaReadBus_req_bits_setIdx,
  input  [18:0] io_metaReadBus_resp_data_0_tag,
  input         io_metaReadBus_resp_data_0_valid,
  input         io_metaReadBus_resp_data_0_dirty,
  input  [18:0] io_metaReadBus_resp_data_1_tag,
  input         io_metaReadBus_resp_data_1_valid,
  input         io_metaReadBus_resp_data_1_dirty,
  input  [18:0] io_metaReadBus_resp_data_2_tag,
  input         io_metaReadBus_resp_data_2_valid,
  input         io_metaReadBus_resp_data_2_dirty,
  input  [18:0] io_metaReadBus_resp_data_3_tag,
  input         io_metaReadBus_resp_data_3_valid,
  input         io_metaReadBus_resp_data_3_dirty,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [9:0]  io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data
);
  wire  _T_29 = io_in_valid & io_metaReadBus_req_ready; // @[Cache.scala 133:31]
  wire  _T_31 = ~io_in_valid; // @[Cache.scala 134:19]
  wire  _T_32 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_33 = _T_31 | _T_32; // @[Cache.scala 134:32]
  wire  _T_34 = _T_33 & io_metaReadBus_req_ready; // @[Cache.scala 134:50]
  assign io_in_ready = _T_34 & io_dataReadBus_req_ready; // @[Cache.scala 134:15]
  assign io_out_valid = _T_29 & io_dataReadBus_req_ready; // @[Cache.scala 133:16]
  assign io_out_bits_req_addr = io_in_bits_addr; // @[Cache.scala 132:19]
  assign io_out_bits_req_size = io_in_bits_size; // @[Cache.scala 132:19]
  assign io_out_bits_req_cmd = io_in_bits_cmd; // @[Cache.scala 132:19]
  assign io_out_bits_req_wmask = io_in_bits_wmask; // @[Cache.scala 132:19]
  assign io_out_bits_req_wdata = io_in_bits_wdata; // @[Cache.scala 132:19]
  assign io_metaReadBus_req_valid = io_in_valid & io_out_ready; // @[SRAMTemplate.scala 53:20]
  assign io_metaReadBus_req_bits_setIdx = io_in_bits_addr[12:6]; // @[SRAMTemplate.scala 26:17]
  assign io_dataReadBus_req_valid = io_in_valid & io_out_ready; // @[SRAMTemplate.scala 53:20]
  assign io_dataReadBus_req_bits_setIdx = {io_in_bits_addr[12:6],io_in_bits_addr[5:3]}; // @[SRAMTemplate.scala 26:17]
endmodule
module CacheStage2_1(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [2:0]  io_in_bits_req_size,
  input  [3:0]  io_in_bits_req_cmd,
  input  [7:0]  io_in_bits_req_wmask,
  input  [63:0] io_in_bits_req_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [2:0]  io_out_bits_req_size,
  output [3:0]  io_out_bits_req_cmd,
  output [7:0]  io_out_bits_req_wmask,
  output [63:0] io_out_bits_req_wdata,
  output [18:0] io_out_bits_metas_0_tag,
  output        io_out_bits_metas_0_valid,
  output        io_out_bits_metas_0_dirty,
  output [18:0] io_out_bits_metas_1_tag,
  output        io_out_bits_metas_1_valid,
  output        io_out_bits_metas_1_dirty,
  output [18:0] io_out_bits_metas_2_tag,
  output        io_out_bits_metas_2_valid,
  output        io_out_bits_metas_2_dirty,
  output [18:0] io_out_bits_metas_3_tag,
  output        io_out_bits_metas_3_valid,
  output        io_out_bits_metas_3_dirty,
  output [63:0] io_out_bits_datas_0_data,
  output [63:0] io_out_bits_datas_1_data,
  output [63:0] io_out_bits_datas_2_data,
  output [63:0] io_out_bits_datas_3_data,
  output        io_out_bits_hit,
  output [3:0]  io_out_bits_waymask,
  output        io_out_bits_mmio,
  output        io_out_bits_isForwardData,
  output [63:0] io_out_bits_forwardData_data_data,
  output [3:0]  io_out_bits_forwardData_waymask,
  input  [18:0] io_metaReadResp_0_tag,
  input         io_metaReadResp_0_valid,
  input         io_metaReadResp_0_dirty,
  input  [18:0] io_metaReadResp_1_tag,
  input         io_metaReadResp_1_valid,
  input         io_metaReadResp_1_dirty,
  input  [18:0] io_metaReadResp_2_tag,
  input         io_metaReadResp_2_valid,
  input         io_metaReadResp_2_dirty,
  input  [18:0] io_metaReadResp_3_tag,
  input         io_metaReadResp_3_valid,
  input         io_metaReadResp_3_dirty,
  input  [63:0] io_dataReadResp_0_data,
  input  [63:0] io_dataReadResp_1_data,
  input  [63:0] io_dataReadResp_2_data,
  input  [63:0] io_dataReadResp_3_data,
  input         io_metaWriteBus_req_valid,
  input  [6:0]  io_metaWriteBus_req_bits_setIdx,
  input  [18:0] io_metaWriteBus_req_bits_data_tag,
  input         io_metaWriteBus_req_bits_data_dirty,
  input  [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_dataWriteBus_req_valid,
  input  [9:0]  io_dataWriteBus_req_bits_setIdx,
  input  [63:0] io_dataWriteBus_req_bits_data_data,
  input  [3:0]  io_dataWriteBus_req_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 162:31]
  wire [6:0] addr_index = io_in_bits_req_addr[12:6]; // @[Cache.scala 162:31]
  wire [18:0] addr_tag = io_in_bits_req_addr[31:13]; // @[Cache.scala 162:31]
  wire  _T_5 = io_in_valid & io_metaWriteBus_req_valid; // @[Cache.scala 164:35]
  wire  _T_12 = io_metaWriteBus_req_bits_setIdx == addr_index; // @[Cache.scala 164:99]
  wire  isForwardMeta = _T_5 & _T_12; // @[Cache.scala 164:64]
  reg  isForwardMetaReg; // @[Cache.scala 165:33]
  wire  _GEN_0 = isForwardMeta | isForwardMetaReg; // @[Cache.scala 166:24]
  wire  _T_13 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire  _T_14 = ~io_in_valid; // @[Cache.scala 167:25]
  wire  _T_15 = _T_13 | _T_14; // @[Cache.scala 167:22]
  reg [18:0] forwardMetaReg_data_tag; // @[Reg.scala 15:16]
  reg  forwardMetaReg_data_dirty; // @[Reg.scala 15:16]
  reg [3:0] forwardMetaReg_waymask; // @[Reg.scala 15:16]
  wire [3:0] _GEN_2 = isForwardMeta ? io_metaWriteBus_req_bits_waymask : forwardMetaReg_waymask; // @[Reg.scala 16:19]
  wire  _GEN_3 = isForwardMeta ? io_metaWriteBus_req_bits_data_dirty : forwardMetaReg_data_dirty; // @[Reg.scala 16:19]
  wire [18:0] _GEN_5 = isForwardMeta ? io_metaWriteBus_req_bits_data_tag : forwardMetaReg_data_tag; // @[Reg.scala 16:19]
  wire  pickForwardMeta = isForwardMetaReg | isForwardMeta; // @[Cache.scala 171:42]
  wire  forwardWaymask_0 = _GEN_2[0]; // @[Cache.scala 173:61]
  wire  forwardWaymask_1 = _GEN_2[1]; // @[Cache.scala 173:61]
  wire  forwardWaymask_2 = _GEN_2[2]; // @[Cache.scala 173:61]
  wire  forwardWaymask_3 = _GEN_2[3]; // @[Cache.scala 173:61]
  wire  _T_16 = pickForwardMeta & forwardWaymask_0; // @[Cache.scala 175:39]
  wire [18:0] metaWay_0_tag = _T_16 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 175:22]
  wire  metaWay_0_valid = _T_16 | io_metaReadResp_0_valid; // @[Cache.scala 175:22]
  wire  _T_18 = pickForwardMeta & forwardWaymask_1; // @[Cache.scala 175:39]
  wire [18:0] metaWay_1_tag = _T_18 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 175:22]
  wire  metaWay_1_valid = _T_18 | io_metaReadResp_1_valid; // @[Cache.scala 175:22]
  wire  _T_20 = pickForwardMeta & forwardWaymask_2; // @[Cache.scala 175:39]
  wire [18:0] metaWay_2_tag = _T_20 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 175:22]
  wire  metaWay_2_valid = _T_20 | io_metaReadResp_2_valid; // @[Cache.scala 175:22]
  wire  _T_22 = pickForwardMeta & forwardWaymask_3; // @[Cache.scala 175:39]
  wire [18:0] metaWay_3_tag = _T_22 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 175:22]
  wire  metaWay_3_valid = _T_22 | io_metaReadResp_3_valid; // @[Cache.scala 175:22]
  wire  _T_24 = metaWay_0_tag == addr_tag; // @[Cache.scala 178:59]
  wire  _T_25 = metaWay_0_valid & _T_24; // @[Cache.scala 178:49]
  wire  _T_26 = _T_25 & io_in_valid; // @[Cache.scala 178:73]
  wire  _T_27 = metaWay_1_tag == addr_tag; // @[Cache.scala 178:59]
  wire  _T_28 = metaWay_1_valid & _T_27; // @[Cache.scala 178:49]
  wire  _T_29 = _T_28 & io_in_valid; // @[Cache.scala 178:73]
  wire  _T_30 = metaWay_2_tag == addr_tag; // @[Cache.scala 178:59]
  wire  _T_31 = metaWay_2_valid & _T_30; // @[Cache.scala 178:49]
  wire  _T_32 = _T_31 & io_in_valid; // @[Cache.scala 178:73]
  wire  _T_33 = metaWay_3_tag == addr_tag; // @[Cache.scala 178:59]
  wire  _T_34 = metaWay_3_valid & _T_33; // @[Cache.scala 178:49]
  wire  _T_35 = _T_34 & io_in_valid; // @[Cache.scala 178:73]
  wire [3:0] hitVec = {_T_35,_T_32,_T_29,_T_26}; // @[Cache.scala 178:90]
  reg [63:0] _T_39; // @[LFSR64.scala 25:23]
  wire  _T_42 = _T_39[0] ^ _T_39[1]; // @[LFSR64.scala 26:23]
  wire  _T_44 = _T_42 ^ _T_39[3]; // @[LFSR64.scala 26:33]
  wire  _T_46 = _T_44 ^ _T_39[4]; // @[LFSR64.scala 26:43]
  wire  _T_47 = _T_39 == 64'h0; // @[LFSR64.scala 28:24]
  wire [63:0] _T_49 = {_T_46,_T_39[63:1]}; // @[Cat.scala 29:58]
  wire [3:0] victimWaymask = 4'h1 << _T_39[1:0]; // @[Cache.scala 179:42]
  wire  _T_52 = ~metaWay_0_valid; // @[Cache.scala 181:45]
  wire  _T_53 = ~metaWay_1_valid; // @[Cache.scala 181:45]
  wire  _T_54 = ~metaWay_2_valid; // @[Cache.scala 181:45]
  wire  _T_55 = ~metaWay_3_valid; // @[Cache.scala 181:45]
  wire [3:0] invalidVec = {_T_55,_T_54,_T_53,_T_52}; // @[Cache.scala 181:56]
  wire  hasInvalidWay = |invalidVec; // @[Cache.scala 182:34]
  wire  _T_59 = invalidVec >= 4'h8; // @[Cache.scala 183:45]
  wire  _T_60 = invalidVec >= 4'h4; // @[Cache.scala 184:20]
  wire  _T_61 = invalidVec >= 4'h2; // @[Cache.scala 185:20]
  wire [1:0] _T_62 = _T_61 ? 2'h2 : 2'h1; // @[Cache.scala 185:8]
  wire [2:0] _T_63 = _T_60 ? 3'h4 : {{1'd0}, _T_62}; // @[Cache.scala 184:8]
  wire [3:0] refillInvalidWaymask = _T_59 ? 4'h8 : {{1'd0}, _T_63}; // @[Cache.scala 183:33]
  wire [3:0] _T_64 = hasInvalidWay ? refillInvalidWaymask : victimWaymask; // @[Cache.scala 188:49]
  wire [3:0] waymask = io_out_bits_hit ? hitVec : _T_64; // @[Cache.scala 188:20]
  wire [1:0] _T_69 = waymask[0] + waymask[1]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_71 = waymask[2] + waymask[3]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_73 = _T_69 + _T_71; // @[Bitwise.scala 47:55]
  wire  _T_75 = _T_73 > 3'h1; // @[Cache.scala 189:26]
  wire  _T_197 = io_in_valid & _T_75; // @[Cache.scala 196:24]
  wire  _T_198 = ~_T_197; // @[Cache.scala 196:10]
  wire  _T_200 = _T_198 | reset; // @[Cache.scala 196:9]
  wire  _T_201 = ~_T_200; // @[Cache.scala 196:9]
  wire  _T_202 = |hitVec; // @[Cache.scala 199:44]
  wire [31:0] _T_204 = io_in_bits_req_addr ^ 32'h30000000; // @[NutCore.scala 86:11]
  wire  _T_206 = _T_204[31:28] == 4'h0; // @[NutCore.scala 86:44]
  wire [31:0] _T_207 = io_in_bits_req_addr ^ 32'he0000000; // @[NutCore.scala 86:11]
  wire  _T_209 = _T_207[31:29] == 3'h0; // @[NutCore.scala 86:44]
  wire [9:0] _T_223 = {addr_index,addr_wordIndex}; // @[Cat.scala 29:58]
  wire  _T_224 = io_dataWriteBus_req_bits_setIdx == _T_223; // @[Cache.scala 205:30]
  wire  _T_225 = io_dataWriteBus_req_valid & _T_224; // @[Cache.scala 205:13]
  wire  isForwardData = io_in_valid & _T_225; // @[Cache.scala 204:35]
  reg  isForwardDataReg; // @[Cache.scala 207:33]
  wire  _GEN_8 = isForwardData | isForwardDataReg; // @[Cache.scala 208:24]
  reg [63:0] forwardDataReg_data_data; // @[Reg.scala 15:16]
  reg [3:0] forwardDataReg_waymask; // @[Reg.scala 15:16]
  wire  _T_232 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign io_in_ready = _T_14 | _T_232; // @[Cache.scala 216:15]
  assign io_out_valid = io_in_valid; // @[Cache.scala 215:16]
  assign io_out_bits_req_addr = io_in_bits_req_addr; // @[Cache.scala 214:19]
  assign io_out_bits_req_size = io_in_bits_req_size; // @[Cache.scala 214:19]
  assign io_out_bits_req_cmd = io_in_bits_req_cmd; // @[Cache.scala 214:19]
  assign io_out_bits_req_wmask = io_in_bits_req_wmask; // @[Cache.scala 214:19]
  assign io_out_bits_req_wdata = io_in_bits_req_wdata; // @[Cache.scala 214:19]
  assign io_out_bits_metas_0_tag = _T_16 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 198:21]
  assign io_out_bits_metas_0_valid = _T_16 | io_metaReadResp_0_valid; // @[Cache.scala 198:21]
  assign io_out_bits_metas_0_dirty = _T_16 ? _GEN_3 : io_metaReadResp_0_dirty; // @[Cache.scala 198:21]
  assign io_out_bits_metas_1_tag = _T_18 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 198:21]
  assign io_out_bits_metas_1_valid = _T_18 | io_metaReadResp_1_valid; // @[Cache.scala 198:21]
  assign io_out_bits_metas_1_dirty = _T_18 ? _GEN_3 : io_metaReadResp_1_dirty; // @[Cache.scala 198:21]
  assign io_out_bits_metas_2_tag = _T_20 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 198:21]
  assign io_out_bits_metas_2_valid = _T_20 | io_metaReadResp_2_valid; // @[Cache.scala 198:21]
  assign io_out_bits_metas_2_dirty = _T_20 ? _GEN_3 : io_metaReadResp_2_dirty; // @[Cache.scala 198:21]
  assign io_out_bits_metas_3_tag = _T_22 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 198:21]
  assign io_out_bits_metas_3_valid = _T_22 | io_metaReadResp_3_valid; // @[Cache.scala 198:21]
  assign io_out_bits_metas_3_dirty = _T_22 ? _GEN_3 : io_metaReadResp_3_dirty; // @[Cache.scala 198:21]
  assign io_out_bits_datas_0_data = io_dataReadResp_0_data; // @[Cache.scala 201:21]
  assign io_out_bits_datas_1_data = io_dataReadResp_1_data; // @[Cache.scala 201:21]
  assign io_out_bits_datas_2_data = io_dataReadResp_2_data; // @[Cache.scala 201:21]
  assign io_out_bits_datas_3_data = io_dataReadResp_3_data; // @[Cache.scala 201:21]
  assign io_out_bits_hit = io_in_valid & _T_202; // @[Cache.scala 199:19]
  assign io_out_bits_waymask = io_out_bits_hit ? hitVec : _T_64; // @[Cache.scala 200:23]
  assign io_out_bits_mmio = _T_206 | _T_209; // @[Cache.scala 202:20]
  assign io_out_bits_isForwardData = isForwardDataReg | isForwardData; // @[Cache.scala 211:29]
  assign io_out_bits_forwardData_data_data = isForwardData ? io_dataWriteBus_req_bits_data_data : forwardDataReg_data_data; // @[Cache.scala 212:27]
  assign io_out_bits_forwardData_waymask = isForwardData ? io_dataWriteBus_req_bits_waymask : forwardDataReg_waymask; // @[Cache.scala 212:27]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  isForwardMetaReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  forwardMetaReg_data_tag = _RAND_1[18:0];
  _RAND_2 = {1{`RANDOM}};
  forwardMetaReg_data_dirty = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  forwardMetaReg_waymask = _RAND_3[3:0];
  _RAND_4 = {2{`RANDOM}};
  _T_39 = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  isForwardDataReg = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  forwardDataReg_data_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  forwardDataReg_waymask = _RAND_7[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      isForwardMetaReg <= 1'h0;
    end else if (_T_15) begin
      isForwardMetaReg <= 1'h0;
    end else begin
      isForwardMetaReg <= _GEN_0;
    end
    if (isForwardMeta) begin
      forwardMetaReg_data_tag <= io_metaWriteBus_req_bits_data_tag;
    end
    if (isForwardMeta) begin
      forwardMetaReg_data_dirty <= io_metaWriteBus_req_bits_data_dirty;
    end
    if (isForwardMeta) begin
      forwardMetaReg_waymask <= io_metaWriteBus_req_bits_waymask;
    end
    if (reset) begin
      _T_39 <= 64'h1234567887654321;
    end else if (_T_47) begin
      _T_39 <= 64'h1;
    end else begin
      _T_39 <= _T_49;
    end
    if (reset) begin
      isForwardDataReg <= 1'h0;
    end else if (_T_15) begin
      isForwardDataReg <= 1'h0;
    end else begin
      isForwardDataReg <= _GEN_8;
    end
    if (isForwardData) begin
      forwardDataReg_data_data <= io_dataWriteBus_req_bits_data_data;
    end
    if (isForwardData) begin
      forwardDataReg_waymask <= io_dataWriteBus_req_bits_waymask;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_201) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Cache.scala:196 assert(!(io.in.valid && PopCount(waymask) > 1.U))\n"); // @[Cache.scala 196:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_201) begin
          $fatal; // @[Cache.scala 196:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CacheStage3_1(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [2:0]  io_in_bits_req_size,
  input  [3:0]  io_in_bits_req_cmd,
  input  [7:0]  io_in_bits_req_wmask,
  input  [63:0] io_in_bits_req_wdata,
  input  [18:0] io_in_bits_metas_0_tag,
  input         io_in_bits_metas_0_valid,
  input         io_in_bits_metas_0_dirty,
  input  [18:0] io_in_bits_metas_1_tag,
  input         io_in_bits_metas_1_valid,
  input         io_in_bits_metas_1_dirty,
  input  [18:0] io_in_bits_metas_2_tag,
  input         io_in_bits_metas_2_valid,
  input         io_in_bits_metas_2_dirty,
  input  [18:0] io_in_bits_metas_3_tag,
  input         io_in_bits_metas_3_valid,
  input         io_in_bits_metas_3_dirty,
  input  [63:0] io_in_bits_datas_0_data,
  input  [63:0] io_in_bits_datas_1_data,
  input  [63:0] io_in_bits_datas_2_data,
  input  [63:0] io_in_bits_datas_3_data,
  input         io_in_bits_hit,
  input  [3:0]  io_in_bits_waymask,
  input         io_in_bits_mmio,
  input         io_in_bits_isForwardData,
  input  [63:0] io_in_bits_forwardData_data_data,
  input  [3:0]  io_in_bits_forwardData_waymask,
  input         io_out_ready,
  output        io_out_valid,
  output [3:0]  io_out_bits_cmd,
  output [63:0] io_out_bits_rdata,
  output        io_isFinish,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [9:0]  io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data,
  output        io_dataWriteBus_req_valid,
  output [9:0]  io_dataWriteBus_req_bits_setIdx,
  output [63:0] io_dataWriteBus_req_bits_data_data,
  output [3:0]  io_dataWriteBus_req_bits_waymask,
  output        io_metaWriteBus_req_valid,
  output [6:0]  io_metaWriteBus_req_bits_setIdx,
  output [18:0] io_metaWriteBus_req_bits_data_tag,
  output        io_metaWriteBus_req_bits_data_dirty,
  output [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [31:0] io_mem_req_bits_addr,
  output [3:0]  io_mem_req_bits_cmd,
  output [63:0] io_mem_req_bits_wdata,
  output        io_mem_resp_ready,
  input         io_mem_resp_valid,
  input  [3:0]  io_mem_resp_bits_cmd,
  input  [63:0] io_mem_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  output [2:0]  io_mmio_req_bits_size,
  output [3:0]  io_mmio_req_bits_cmd,
  output [7:0]  io_mmio_req_bits_wmask,
  output [63:0] io_mmio_req_bits_wdata,
  output        io_mmio_resp_ready,
  input         io_mmio_resp_valid,
  input  [63:0] io_mmio_resp_bits_rdata,
  output        io_cohResp_valid,
  output [3:0]  io_cohResp_bits_cmd,
  output [63:0] io_cohResp_bits_rdata,
  output        io_dataReadRespToL1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  metaWriteArb_io_in_0_valid; // @[Cache.scala 241:28]
  wire [6:0] metaWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 241:28]
  wire [18:0] metaWriteArb_io_in_0_bits_data_tag; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_in_0_bits_data_dirty; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_in_0_bits_waymask; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_in_1_valid; // @[Cache.scala 241:28]
  wire [6:0] metaWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 241:28]
  wire [18:0] metaWriteArb_io_in_1_bits_data_tag; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_in_1_bits_data_dirty; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_in_1_bits_waymask; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_out_valid; // @[Cache.scala 241:28]
  wire [6:0] metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 241:28]
  wire [18:0] metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_out_bits_waymask; // @[Cache.scala 241:28]
  wire  dataWriteArb_io_in_0_valid; // @[Cache.scala 242:28]
  wire [9:0] dataWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 242:28]
  wire [63:0] dataWriteArb_io_in_0_bits_data_data; // @[Cache.scala 242:28]
  wire [3:0] dataWriteArb_io_in_0_bits_waymask; // @[Cache.scala 242:28]
  wire  dataWriteArb_io_in_1_valid; // @[Cache.scala 242:28]
  wire [9:0] dataWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 242:28]
  wire [63:0] dataWriteArb_io_in_1_bits_data_data; // @[Cache.scala 242:28]
  wire [3:0] dataWriteArb_io_in_1_bits_waymask; // @[Cache.scala 242:28]
  wire  dataWriteArb_io_out_valid; // @[Cache.scala 242:28]
  wire [9:0] dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 242:28]
  wire [63:0] dataWriteArb_io_out_bits_data_data; // @[Cache.scala 242:28]
  wire [3:0] dataWriteArb_io_out_bits_waymask; // @[Cache.scala 242:28]
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 245:31]
  wire [6:0] addr_index = io_in_bits_req_addr[12:6]; // @[Cache.scala 245:31]
  wire  mmio = io_in_valid & io_in_bits_mmio; // @[Cache.scala 246:26]
  wire  hit = io_in_valid & io_in_bits_hit; // @[Cache.scala 247:25]
  wire  _T_5 = ~io_in_bits_hit; // @[Cache.scala 248:29]
  wire  miss = io_in_valid & _T_5; // @[Cache.scala 248:26]
  wire  _T_7 = io_in_bits_req_cmd == 4'h8; // @[SimpleBus.scala 79:23]
  wire  probe = io_in_valid & _T_7; // @[Cache.scala 249:39]
  wire  _T_8 = io_in_bits_req_cmd == 4'h2; // @[SimpleBus.scala 76:27]
  wire  hitReadBurst = hit & _T_8; // @[Cache.scala 250:26]
  wire [20:0] _T_14 = {io_in_bits_metas_0_tag,io_in_bits_metas_0_valid,io_in_bits_metas_0_dirty}; // @[Mux.scala 27:72]
  wire [20:0] _T_15 = io_in_bits_waymask[0] ? _T_14 : 21'h0; // @[Mux.scala 27:72]
  wire [20:0] _T_17 = {io_in_bits_metas_1_tag,io_in_bits_metas_1_valid,io_in_bits_metas_1_dirty}; // @[Mux.scala 27:72]
  wire [20:0] _T_18 = io_in_bits_waymask[1] ? _T_17 : 21'h0; // @[Mux.scala 27:72]
  wire [20:0] _T_20 = {io_in_bits_metas_2_tag,io_in_bits_metas_2_valid,io_in_bits_metas_2_dirty}; // @[Mux.scala 27:72]
  wire [20:0] _T_21 = io_in_bits_waymask[2] ? _T_20 : 21'h0; // @[Mux.scala 27:72]
  wire [20:0] _T_23 = {io_in_bits_metas_3_tag,io_in_bits_metas_3_valid,io_in_bits_metas_3_dirty}; // @[Mux.scala 27:72]
  wire [20:0] _T_24 = io_in_bits_waymask[3] ? _T_23 : 21'h0; // @[Mux.scala 27:72]
  wire [20:0] _T_25 = _T_15 | _T_18; // @[Mux.scala 27:72]
  wire [20:0] _T_26 = _T_25 | _T_21; // @[Mux.scala 27:72]
  wire [20:0] _T_27 = _T_26 | _T_24; // @[Mux.scala 27:72]
  wire  meta_dirty = _T_27[0]; // @[Mux.scala 27:72]
  wire [18:0] meta_tag = _T_27[20:2]; // @[Mux.scala 27:72]
  wire  _T_32 = mmio & hit; // @[Cache.scala 252:17]
  wire  _T_33 = ~_T_32; // @[Cache.scala 252:10]
  wire  _T_35 = _T_33 | reset; // @[Cache.scala 252:9]
  wire  _T_36 = ~_T_35; // @[Cache.scala 252:9]
  wire  _T_37 = io_in_bits_waymask == io_in_bits_forwardData_waymask; // @[Cache.scala 260:71]
  wire  useForwardData = io_in_bits_isForwardData & _T_37; // @[Cache.scala 260:49]
  wire [63:0] _T_42 = io_in_bits_waymask[0] ? io_in_bits_datas_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_43 = io_in_bits_waymask[1] ? io_in_bits_datas_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_44 = io_in_bits_waymask[2] ? io_in_bits_datas_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_45 = io_in_bits_waymask[3] ? io_in_bits_datas_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_46 = _T_42 | _T_43; // @[Mux.scala 27:72]
  wire [63:0] _T_47 = _T_46 | _T_44; // @[Mux.scala 27:72]
  wire [63:0] _T_48 = _T_47 | _T_45; // @[Mux.scala 27:72]
  wire [63:0] dataRead = useForwardData ? io_in_bits_forwardData_data_data : _T_48; // @[Cache.scala 262:21]
  wire [7:0] _T_64 = io_in_bits_req_wmask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_66 = io_in_bits_req_wmask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_68 = io_in_bits_req_wmask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_70 = io_in_bits_req_wmask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_72 = io_in_bits_req_wmask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_74 = io_in_bits_req_wmask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_76 = io_in_bits_req_wmask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_78 = io_in_bits_req_wmask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_85 = {_T_78,_T_76,_T_74,_T_72,_T_70,_T_68,_T_66,_T_64}; // @[Cat.scala 29:58]
  wire [63:0] wordMask = io_in_bits_req_cmd[0] ? _T_85 : 64'h0; // @[Cache.scala 263:21]
  reg [2:0] value; // @[Counter.scala 29:33]
  wire  _T_86 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_87 = io_in_bits_req_cmd == 4'h3; // @[Cache.scala 266:34]
  wire  _T_88 = io_in_bits_req_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_89 = _T_87 | _T_88; // @[Cache.scala 266:62]
  wire  _T_90 = _T_86 & _T_89; // @[Cache.scala 266:22]
  wire [2:0] _T_93 = value + 3'h1; // @[Counter.scala 39:22]
  wire [2:0] _GEN_0 = _T_90 ? _T_93 : value; // @[Cache.scala 266:85]
  wire  hitWrite = hit & io_in_bits_req_cmd[0]; // @[Cache.scala 270:22]
  wire [63:0] _T_96 = io_in_bits_req_wdata & wordMask; // @[BitUtils.scala 32:13]
  wire [63:0] _T_97 = ~wordMask; // @[BitUtils.scala 32:38]
  wire [63:0] _T_98 = dataRead & _T_97; // @[BitUtils.scala 32:36]
  wire [2:0] _T_103 = _T_89 ? value : addr_wordIndex; // @[Cache.scala 273:51]
  wire  _T_105 = ~meta_dirty; // @[Cache.scala 276:25]
  wire  metaHitWriteBus_req_valid = hitWrite & _T_105; // @[Cache.scala 276:22]
  reg [3:0] state; // @[Cache.scala 281:22]
  reg [2:0] value_1; // @[Counter.scala 29:33]
  reg [2:0] value_2; // @[Counter.scala 29:33]
  reg [1:0] state2; // @[Cache.scala 291:23]
  wire  _T_118 = state == 4'h3; // @[Cache.scala 293:39]
  wire  _T_119 = state == 4'h8; // @[Cache.scala 293:66]
  wire  _T_120 = _T_118 | _T_119; // @[Cache.scala 293:57]
  wire  _T_121 = state2 == 2'h0; // @[Cache.scala 293:92]
  wire [2:0] _T_124 = _T_119 ? value_1 : value_2; // @[Cache.scala 294:33]
  wire  _T_126 = state2 == 2'h1; // @[Cache.scala 295:60]
  reg [63:0] dataWay_0_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_1_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_2_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_3_data; // @[Reg.scala 15:16]
  wire [63:0] _T_131 = io_in_bits_waymask[0] ? dataWay_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_132 = io_in_bits_waymask[1] ? dataWay_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_133 = io_in_bits_waymask[2] ? dataWay_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_134 = io_in_bits_waymask[3] ? dataWay_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_135 = _T_131 | _T_132; // @[Mux.scala 27:72]
  wire [63:0] _T_136 = _T_135 | _T_133; // @[Mux.scala 27:72]
  wire  _T_141 = 2'h0 == state2; // @[Conditional.scala 37:30]
  wire  _T_142 = io_dataReadBus_req_ready & io_dataReadBus_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_143 = 2'h1 == state2; // @[Conditional.scala 37:30]
  wire  _T_144 = 2'h2 == state2; // @[Conditional.scala 37:30]
  wire  _T_145 = io_mem_req_ready & io_mem_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_147 = _T_145 | io_cohResp_valid; // @[Cache.scala 301:46]
  wire  _T_148 = hitReadBurst & io_out_ready; // @[Cache.scala 301:83]
  wire  _T_149 = _T_147 | _T_148; // @[Cache.scala 301:67]
  wire [31:0] raddr = {io_in_bits_req_addr[31:3],3'h0}; // @[Cat.scala 29:58]
  wire [31:0] waddr = {meta_tag,addr_index,6'h0}; // @[Cat.scala 29:58]
  wire  _T_152 = state == 4'h1; // @[Cache.scala 309:23]
  wire  _T_153 = value_2 == 3'h7; // @[Cache.scala 310:29]
  wire [2:0] _T_154 = _T_153 ? 3'h7 : 3'h3; // @[Cache.scala 310:8]
  wire [2:0] cmd = _T_152 ? 3'h2 : _T_154; // @[Cache.scala 309:16]
  wire  _T_160 = state2 == 2'h2; // @[Cache.scala 316:89]
  wire  _T_161 = _T_118 & _T_160; // @[Cache.scala 316:78]
  reg  afterFirstRead; // @[Cache.scala 323:31]
  reg  alreadyOutFire; // @[Reg.scala 27:20]
  wire  _GEN_12 = _T_86 | alreadyOutFire; // @[Reg.scala 28:19]
  wire  _T_165 = ~afterFirstRead; // @[Cache.scala 325:22]
  wire  _T_166 = io_mem_resp_ready & io_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_167 = _T_165 & _T_166; // @[Cache.scala 325:38]
  wire  _T_168 = state == 4'h2; // @[Cache.scala 325:70]
  wire  readingFirst = _T_167 & _T_168; // @[Cache.scala 325:60]
  wire  _T_170 = state == 4'h6; // @[Cache.scala 327:52]
  wire  _T_171 = mmio ? _T_170 : readingFirst; // @[Cache.scala 327:39]
  reg [63:0] inRdataRegDemand; // @[Reg.scala 15:16]
  wire  _T_172 = state == 4'h0; // @[Cache.scala 330:31]
  wire  _T_173 = _T_172 & probe; // @[Cache.scala 330:43]
  wire  _T_176 = _T_119 & _T_160; // @[Cache.scala 331:46]
  wire  _T_180 = _T_119 & io_cohResp_valid; // @[Cache.scala 333:49]
  reg [2:0] _T_181; // @[Counter.scala 29:33]
  wire  _T_182 = _T_181 == 3'h7; // @[Counter.scala 38:24]
  wire [2:0] _T_184 = _T_181 + 3'h1; // @[Counter.scala 39:22]
  wire  releaseLast = _T_180 & _T_182; // @[Counter.scala 67:17]
  wire [2:0] _T_186 = releaseLast ? 3'h6 : 3'h0; // @[Cache.scala 334:54]
  wire [3:0] _T_187 = hit ? 4'hc : 4'h8; // @[Cache.scala 335:8]
  wire  respToL1Fire = _T_148 & _T_160; // @[Cache.scala 337:51]
  wire  _T_195 = _T_172 | _T_176; // @[Cache.scala 338:48]
  wire  _T_196 = _T_195 & hitReadBurst; // @[Cache.scala 338:96]
  wire  _T_197 = _T_196 & io_out_ready; // @[Cache.scala 338:112]
  reg [2:0] _T_198; // @[Counter.scala 29:33]
  wire  _T_199 = _T_198 == 3'h7; // @[Counter.scala 38:24]
  wire [2:0] _T_201 = _T_198 + 3'h1; // @[Counter.scala 39:22]
  wire  respToL1Last = _T_197 & _T_199; // @[Counter.scala 67:17]
  wire  _T_202 = 4'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_206 = addr_wordIndex == 3'h7; // @[Cache.scala 352:49]
  wire [2:0] _T_208 = addr_wordIndex + 3'h1; // @[Cache.scala 352:93]
  wire  _T_210 = miss | mmio; // @[Cache.scala 353:26]
  wire  _T_217 = 4'h5 == state; // @[Conditional.scala 37:30]
  wire  _T_218 = io_mmio_req_ready & io_mmio_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_219 = 4'h6 == state; // @[Conditional.scala 37:30]
  wire  _T_220 = io_mmio_resp_ready & io_mmio_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_221 = 4'h8 == state; // @[Conditional.scala 37:30]
  wire  _T_223 = io_cohResp_valid | respToL1Fire; // @[Cache.scala 362:31]
  wire [2:0] _T_226 = value_1 + 3'h1; // @[Counter.scala 39:22]
  wire  _T_228 = probe & io_cohResp_valid; // @[Cache.scala 363:19]
  wire  _T_229 = _T_228 & releaseLast; // @[Cache.scala 363:40]
  wire  _T_230 = respToL1Fire & respToL1Last; // @[Cache.scala 363:71]
  wire  _T_231 = _T_229 | _T_230; // @[Cache.scala 363:55]
  wire  _T_232 = 4'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_234 = 4'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_240 = io_mem_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire  _GEN_33 = _T_166 | afterFirstRead; // @[Cache.scala 372:33]
  wire  _T_241 = 4'h3 == state; // @[Conditional.scala 37:30]
  wire [2:0] _T_245 = value_2 + 3'h1; // @[Counter.scala 39:22]
  wire  _T_246 = io_mem_req_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_248 = _T_246 & _T_145; // @[Cache.scala 382:43]
  wire  _T_249 = 4'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_251 = 4'h7 == state; // @[Conditional.scala 37:30]
  wire [63:0] _T_255 = readingFirst ? wordMask : 64'h0; // @[Cache.scala 389:67]
  wire [63:0] _T_256 = io_in_bits_req_wdata & _T_255; // @[BitUtils.scala 32:13]
  wire [63:0] _T_257 = ~_T_255; // @[BitUtils.scala 32:38]
  wire [63:0] _T_258 = io_mem_resp_bits_rdata & _T_257; // @[BitUtils.scala 32:36]
  wire  dataRefillWriteBus_req_valid = _T_168 & _T_166; // @[Cache.scala 391:39]
  wire  metaRefillWriteBus_req_valid = dataRefillWriteBus_req_valid & _T_240; // @[Cache.scala 399:61]
  wire  _T_281 = ~io_in_bits_req_cmd[0]; // @[SimpleBus.scala 73:18]
  wire  _T_283 = ~io_in_bits_req_cmd[3]; // @[SimpleBus.scala 73:29]
  wire  _T_284 = _T_281 & _T_283; // @[SimpleBus.scala 73:26]
  wire [2:0] _T_286 = io_in_bits_req_cmd[0] ? 3'h5 : 3'h0; // @[Cache.scala 427:79]
  wire [2:0] _T_288 = _T_284 ? 3'h6 : _T_286; // @[Cache.scala 427:27]
  wire  _T_293 = state == 4'h7; // @[Cache.scala 433:48]
  wire  _T_308 = io_in_bits_req_cmd[0] | mmio; // @[Cache.scala 434:60]
  wire  _T_310 = ~alreadyOutFire; // @[Cache.scala 434:110]
  wire  _T_311 = afterFirstRead & _T_310; // @[Cache.scala 434:107]
  wire  _T_312 = _T_308 ? _T_293 : _T_311; // @[Cache.scala 434:45]
  wire  _T_313 = hit | _T_312; // @[Cache.scala 434:28]
  wire  _T_314 = probe ? 1'h0 : _T_313; // @[Cache.scala 434:8]
  wire  _T_320 = _T_119 & releaseLast; // @[Cache.scala 441:100]
  wire  _T_321 = miss ? _T_172 : _T_320; // @[Cache.scala 441:53]
  wire  _T_322 = io_cohResp_valid & _T_321; // @[Cache.scala 441:47]
  wire  _T_324 = hit | io_in_bits_req_cmd[0]; // @[Cache.scala 442:13]
  wire  _T_329 = _T_293 & _GEN_12; // @[Cache.scala 442:70]
  wire  _T_330 = _T_324 ? _T_86 : _T_329; // @[Cache.scala 442:8]
  wire  _T_333 = ~hitReadBurst; // @[Cache.scala 445:55]
  wire  _T_334 = _T_172 & _T_333; // @[Cache.scala 445:52]
  wire  _T_335 = io_out_ready & _T_334; // @[Cache.scala 445:31]
  wire  _T_336 = ~miss; // @[Cache.scala 445:73]
  wire  _T_337 = _T_335 & _T_336; // @[Cache.scala 445:70]
  wire  _T_338 = ~probe; // @[Cache.scala 445:82]
  wire  _T_341 = _T_172 & io_out_ready; // @[Cache.scala 446:60]
  wire  _T_345 = _T_341 | _T_176; // @[Cache.scala 446:76]
  wire  _T_347 = metaHitWriteBus_req_valid & metaRefillWriteBus_req_valid; // @[Cache.scala 448:38]
  wire  _T_348 = ~_T_347; // @[Cache.scala 448:10]
  wire  _T_350 = _T_348 | reset; // @[Cache.scala 448:9]
  wire  _T_351 = ~_T_350; // @[Cache.scala 448:9]
  wire  _T_352 = hitWrite & dataRefillWriteBus_req_valid; // @[Cache.scala 449:38]
  wire  _T_353 = ~_T_352; // @[Cache.scala 449:10]
  wire  _T_355 = _T_353 | reset; // @[Cache.scala 449:9]
  wire  _T_356 = ~_T_355; // @[Cache.scala 449:9]
  Arbiter metaWriteArb ( // @[Cache.scala 241:28]
    .io_in_0_valid(metaWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(metaWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_tag(metaWriteArb_io_in_0_bits_data_tag),
    .io_in_0_bits_data_dirty(metaWriteArb_io_in_0_bits_data_dirty),
    .io_in_0_bits_waymask(metaWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(metaWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(metaWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_tag(metaWriteArb_io_in_1_bits_data_tag),
    .io_in_1_bits_data_dirty(metaWriteArb_io_in_1_bits_data_dirty),
    .io_in_1_bits_waymask(metaWriteArb_io_in_1_bits_waymask),
    .io_out_valid(metaWriteArb_io_out_valid),
    .io_out_bits_setIdx(metaWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_tag(metaWriteArb_io_out_bits_data_tag),
    .io_out_bits_data_dirty(metaWriteArb_io_out_bits_data_dirty),
    .io_out_bits_waymask(metaWriteArb_io_out_bits_waymask)
  );
  Arbiter_1 dataWriteArb ( // @[Cache.scala 242:28]
    .io_in_0_valid(dataWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(dataWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_data(dataWriteArb_io_in_0_bits_data_data),
    .io_in_0_bits_waymask(dataWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(dataWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(dataWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_data(dataWriteArb_io_in_1_bits_data_data),
    .io_in_1_bits_waymask(dataWriteArb_io_in_1_bits_waymask),
    .io_out_valid(dataWriteArb_io_out_valid),
    .io_out_bits_setIdx(dataWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_data(dataWriteArb_io_out_bits_data_data),
    .io_out_bits_waymask(dataWriteArb_io_out_bits_waymask)
  );
  assign io_in_ready = _T_337 & _T_338; // @[Cache.scala 445:15]
  assign io_out_valid = io_in_valid & _T_314; // @[Cache.scala 432:16]
  assign io_out_bits_cmd = {{1'd0}, _T_288}; // @[Cache.scala 427:21]
  assign io_out_bits_rdata = hit ? dataRead : inRdataRegDemand; // @[Cache.scala 426:23]
  assign io_isFinish = probe ? _T_322 : _T_330; // @[Cache.scala 441:15]
  assign io_dataReadBus_req_valid = _T_120 & _T_121; // @[SRAMTemplate.scala 53:20]
  assign io_dataReadBus_req_bits_setIdx = {addr_index,_T_124}; // @[SRAMTemplate.scala 26:17]
  assign io_dataWriteBus_req_valid = dataWriteArb_io_out_valid; // @[Cache.scala 396:23]
  assign io_dataWriteBus_req_bits_setIdx = dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 396:23]
  assign io_dataWriteBus_req_bits_data_data = dataWriteArb_io_out_bits_data_data; // @[Cache.scala 396:23]
  assign io_dataWriteBus_req_bits_waymask = dataWriteArb_io_out_bits_waymask; // @[Cache.scala 396:23]
  assign io_metaWriteBus_req_valid = metaWriteArb_io_out_valid; // @[Cache.scala 406:23]
  assign io_metaWriteBus_req_bits_setIdx = metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 406:23]
  assign io_metaWriteBus_req_bits_data_tag = metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 406:23]
  assign io_metaWriteBus_req_bits_data_dirty = metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 406:23]
  assign io_metaWriteBus_req_bits_waymask = metaWriteArb_io_out_bits_waymask; // @[Cache.scala 406:23]
  assign io_mem_req_valid = _T_152 | _T_161; // @[Cache.scala 316:20]
  assign io_mem_req_bits_addr = _T_152 ? raddr : waddr; // @[SimpleBus.scala 64:15]
  assign io_mem_req_bits_cmd = {{1'd0}, cmd}; // @[SimpleBus.scala 65:14]
  assign io_mem_req_bits_wdata = _T_136 | _T_134; // @[SimpleBus.scala 67:16]
  assign io_mem_resp_ready = 1'h1; // @[Cache.scala 315:21]
  assign io_mmio_req_valid = state == 4'h5; // @[Cache.scala 321:21]
  assign io_mmio_req_bits_addr = io_in_bits_req_addr; // @[Cache.scala 319:20]
  assign io_mmio_req_bits_size = io_in_bits_req_size; // @[Cache.scala 319:20]
  assign io_mmio_req_bits_cmd = io_in_bits_req_cmd; // @[Cache.scala 319:20]
  assign io_mmio_req_bits_wmask = io_in_bits_req_wmask; // @[Cache.scala 319:20]
  assign io_mmio_req_bits_wdata = io_in_bits_req_wdata; // @[Cache.scala 319:20]
  assign io_mmio_resp_ready = 1'h1; // @[Cache.scala 320:22]
  assign io_cohResp_valid = _T_173 | _T_176; // @[Cache.scala 330:20]
  assign io_cohResp_bits_cmd = _T_119 ? {{1'd0}, _T_186} : _T_187; // @[Cache.scala 334:23]
  assign io_cohResp_bits_rdata = _T_136 | _T_134; // @[Cache.scala 332:25]
  assign io_dataReadRespToL1 = hitReadBurst & _T_345; // @[Cache.scala 446:23]
  assign metaWriteArb_io_in_0_valid = hitWrite & _T_105; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_0_bits_setIdx = io_in_bits_req_addr[12:6]; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_0_bits_data_tag = _T_27[20:2]; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_0_bits_data_dirty = 1'h1; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_1_valid = dataRefillWriteBus_req_valid & _T_240; // @[Cache.scala 405:25]
  assign metaWriteArb_io_in_1_bits_setIdx = io_in_bits_req_addr[12:6]; // @[Cache.scala 405:25]
  assign metaWriteArb_io_in_1_bits_data_tag = io_in_bits_req_addr[31:13]; // @[Cache.scala 405:25]
  assign metaWriteArb_io_in_1_bits_data_dirty = io_in_bits_req_cmd[0]; // @[Cache.scala 405:25]
  assign metaWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 405:25]
  assign dataWriteArb_io_in_0_valid = hit & io_in_bits_req_cmd[0]; // @[Cache.scala 394:25]
  assign dataWriteArb_io_in_0_bits_setIdx = {addr_index,_T_103}; // @[Cache.scala 394:25]
  assign dataWriteArb_io_in_0_bits_data_data = _T_96 | _T_98; // @[Cache.scala 394:25]
  assign dataWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 394:25]
  assign dataWriteArb_io_in_1_valid = _T_168 & _T_166; // @[Cache.scala 395:25]
  assign dataWriteArb_io_in_1_bits_setIdx = {addr_index,value_1}; // @[Cache.scala 395:25]
  assign dataWriteArb_io_in_1_bits_data_data = _T_256 | _T_258; // @[Cache.scala 395:25]
  assign dataWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 395:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  value_2 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  state2 = _RAND_4[1:0];
  _RAND_5 = {2{`RANDOM}};
  dataWay_0_data = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  dataWay_1_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  dataWay_2_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  dataWay_3_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  afterFirstRead = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  alreadyOutFire = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  inRdataRegDemand = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  _T_181 = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  _T_198 = _RAND_13[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 3'h0;
    end else if (_T_202) begin
      if (_T_90) begin
        value <= _T_93;
      end
    end else if (_T_217) begin
      if (_T_90) begin
        value <= _T_93;
      end
    end else if (_T_219) begin
      if (_T_90) begin
        value <= _T_93;
      end
    end else if (_T_221) begin
      if (_T_90) begin
        value <= _T_93;
      end
    end else if (_T_232) begin
      value <= _GEN_0;
    end else if (_T_234) begin
      if (_T_166) begin
        if (_T_87) begin
          value <= 3'h0;
        end else begin
          value <= _GEN_0;
        end
      end else begin
        value <= _GEN_0;
      end
    end else begin
      value <= _GEN_0;
    end
    if (reset) begin
      state <= 4'h0;
    end else if (_T_202) begin
      if (probe) begin
        if (io_cohResp_valid) begin
          if (hit) begin
            state <= 4'h8;
          end else begin
            state <= 4'h0;
          end
        end
      end else if (_T_148) begin
        state <= 4'h8;
      end else if (_T_210) begin
        if (mmio) begin
          state <= 4'h5;
        end else if (meta_dirty) begin
          state <= 4'h3;
        end else begin
          state <= 4'h1;
        end
      end
    end else if (_T_217) begin
      if (_T_218) begin
        state <= 4'h6;
      end
    end else if (_T_219) begin
      if (_T_220) begin
        state <= 4'h7;
      end
    end else if (_T_221) begin
      if (_T_231) begin
        state <= 4'h0;
      end
    end else if (_T_232) begin
      if (_T_145) begin
        state <= 4'h2;
      end
    end else if (_T_234) begin
      if (_T_166) begin
        if (_T_240) begin
          state <= 4'h7;
        end
      end
    end else if (_T_241) begin
      if (_T_248) begin
        state <= 4'h4;
      end
    end else if (_T_249) begin
      if (_T_166) begin
        state <= 4'h1;
      end
    end else if (_T_251) begin
      if (_GEN_12) begin
        state <= 4'h0;
      end
    end
    if (reset) begin
      value_1 <= 3'h0;
    end else if (_T_202) begin
      if (probe) begin
        if (io_cohResp_valid) begin
          value_1 <= addr_wordIndex;
        end
      end else if (_T_148) begin
        if (_T_206) begin
          value_1 <= 3'h0;
        end else begin
          value_1 <= _T_208;
        end
      end
    end else if (!(_T_217)) begin
      if (!(_T_219)) begin
        if (_T_221) begin
          if (_T_223) begin
            value_1 <= _T_226;
          end
        end else if (_T_232) begin
          if (_T_145) begin
            value_1 <= addr_wordIndex;
          end
        end else if (_T_234) begin
          if (_T_166) begin
            value_1 <= _T_226;
          end
        end
      end
    end
    if (reset) begin
      value_2 <= 3'h0;
    end else if (!(_T_202)) begin
      if (!(_T_217)) begin
        if (!(_T_219)) begin
          if (!(_T_221)) begin
            if (!(_T_232)) begin
              if (!(_T_234)) begin
                if (_T_241) begin
                  if (_T_145) begin
                    value_2 <= _T_245;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      state2 <= 2'h0;
    end else if (_T_141) begin
      if (_T_142) begin
        state2 <= 2'h1;
      end
    end else if (_T_143) begin
      state2 <= 2'h2;
    end else if (_T_144) begin
      if (_T_149) begin
        state2 <= 2'h0;
      end
    end
    if (_T_126) begin
      dataWay_0_data <= io_dataReadBus_resp_data_0_data;
    end
    if (_T_126) begin
      dataWay_1_data <= io_dataReadBus_resp_data_1_data;
    end
    if (_T_126) begin
      dataWay_2_data <= io_dataReadBus_resp_data_2_data;
    end
    if (_T_126) begin
      dataWay_3_data <= io_dataReadBus_resp_data_3_data;
    end
    if (reset) begin
      afterFirstRead <= 1'h0;
    end else if (_T_202) begin
      afterFirstRead <= 1'h0;
    end else if (!(_T_217)) begin
      if (!(_T_219)) begin
        if (!(_T_221)) begin
          if (!(_T_232)) begin
            if (_T_234) begin
              afterFirstRead <= _GEN_33;
            end
          end
        end
      end
    end
    if (reset) begin
      alreadyOutFire <= 1'h0;
    end else if (_T_202) begin
      alreadyOutFire <= 1'h0;
    end else begin
      alreadyOutFire <= _GEN_12;
    end
    if (_T_171) begin
      if (mmio) begin
        inRdataRegDemand <= io_mmio_resp_bits_rdata;
      end else begin
        inRdataRegDemand <= io_mem_resp_bits_rdata;
      end
    end
    if (reset) begin
      _T_181 <= 3'h0;
    end else if (_T_180) begin
      _T_181 <= _T_184;
    end
    if (reset) begin
      _T_198 <= 3'h0;
    end else if (_T_197) begin
      _T_198 <= _T_201;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_36) begin
          $fwrite(32'h80000002,"Assertion failed: MMIO request should not hit in cache\n    at Cache.scala:252 assert(!(mmio && hit), \"MMIO request should not hit in cache\")\n"); // @[Cache.scala 252:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_36) begin
          $fatal; // @[Cache.scala 252:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_351) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Cache.scala:448 assert(!(metaHitWriteBus.req.valid && metaRefillWriteBus.req.valid))\n"); // @[Cache.scala 448:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_351) begin
          $fatal; // @[Cache.scala 448:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_356) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Cache.scala:449 assert(!(dataHitWriteBus.req.valid && dataRefillWriteBus.req.valid))\n"); // @[Cache.scala 449:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_356) begin
          $fatal; // @[Cache.scala 449:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Arbiter_9(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [31:0] io_in_0_bits_addr,
  input  [2:0]  io_in_0_bits_size,
  input  [3:0]  io_in_0_bits_cmd,
  input  [7:0]  io_in_0_bits_wmask,
  input  [63:0] io_in_0_bits_wdata,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [31:0] io_in_1_bits_addr,
  input  [2:0]  io_in_1_bits_size,
  input  [3:0]  io_in_1_bits_cmd,
  input  [7:0]  io_in_1_bits_wmask,
  input  [63:0] io_in_1_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [2:0]  io_out_bits_size,
  output [3:0]  io_out_bits_cmd,
  output [7:0]  io_out_bits_wmask,
  output [63:0] io_out_bits_wdata
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  _T_2 = ~grant_1; // @[Arbiter.scala 135:19]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = _T_2 | io_in_1_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_addr = io_in_0_valid ? io_in_0_bits_addr : io_in_1_bits_addr; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_size = io_in_0_valid ? io_in_0_bits_size : io_in_1_bits_size; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_cmd = io_in_0_valid ? io_in_0_bits_cmd : io_in_1_bits_cmd; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_wmask = io_in_0_valid ? io_in_0_bits_wmask : io_in_1_bits_wmask; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_wdata = io_in_0_valid ? io_in_0_bits_wdata : io_in_1_bits_wdata; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
endmodule
module Cache_1(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_mem_req_ready,
  output        io_out_mem_req_valid,
  output [31:0] io_out_mem_req_bits_addr,
  output [3:0]  io_out_mem_req_bits_cmd,
  output [63:0] io_out_mem_req_bits_wdata,
  input         io_out_mem_resp_valid,
  input  [3:0]  io_out_mem_resp_bits_cmd,
  input  [63:0] io_out_mem_resp_bits_rdata,
  output        io_out_coh_req_ready,
  input         io_out_coh_req_valid,
  input  [31:0] io_out_coh_req_bits_addr,
  input  [63:0] io_out_coh_req_bits_wdata,
  output        io_out_coh_resp_valid,
  output [3:0]  io_out_coh_resp_bits_cmd,
  output [63:0] io_out_coh_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  output [2:0]  io_mmio_req_bits_size,
  output [3:0]  io_mmio_req_bits_cmd,
  output [7:0]  io_mmio_req_bits_wmask,
  output [63:0] io_mmio_req_bits_wdata,
  input         io_mmio_resp_valid,
  input  [63:0] io_mmio_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [63:0] _RAND_26;
  reg [63:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [31:0] _RAND_30;
  reg [31:0] _RAND_31;
  reg [63:0] _RAND_32;
  reg [31:0] _RAND_33;
`endif // RANDOMIZE_REG_INIT
  wire  s1_io_in_ready; // @[Cache.scala 475:18]
  wire  s1_io_in_valid; // @[Cache.scala 475:18]
  wire [31:0] s1_io_in_bits_addr; // @[Cache.scala 475:18]
  wire [2:0] s1_io_in_bits_size; // @[Cache.scala 475:18]
  wire [3:0] s1_io_in_bits_cmd; // @[Cache.scala 475:18]
  wire [7:0] s1_io_in_bits_wmask; // @[Cache.scala 475:18]
  wire [63:0] s1_io_in_bits_wdata; // @[Cache.scala 475:18]
  wire  s1_io_out_ready; // @[Cache.scala 475:18]
  wire  s1_io_out_valid; // @[Cache.scala 475:18]
  wire [31:0] s1_io_out_bits_req_addr; // @[Cache.scala 475:18]
  wire [2:0] s1_io_out_bits_req_size; // @[Cache.scala 475:18]
  wire [3:0] s1_io_out_bits_req_cmd; // @[Cache.scala 475:18]
  wire [7:0] s1_io_out_bits_req_wmask; // @[Cache.scala 475:18]
  wire [63:0] s1_io_out_bits_req_wdata; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_req_ready; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_req_valid; // @[Cache.scala 475:18]
  wire [6:0] s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 475:18]
  wire [18:0] s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_0_dirty; // @[Cache.scala 475:18]
  wire [18:0] s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_1_dirty; // @[Cache.scala 475:18]
  wire [18:0] s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_2_dirty; // @[Cache.scala 475:18]
  wire [18:0] s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_3_dirty; // @[Cache.scala 475:18]
  wire  s1_io_dataReadBus_req_ready; // @[Cache.scala 475:18]
  wire  s1_io_dataReadBus_req_valid; // @[Cache.scala 475:18]
  wire [9:0] s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 475:18]
  wire [63:0] s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 475:18]
  wire [63:0] s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 475:18]
  wire [63:0] s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 475:18]
  wire [63:0] s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 475:18]
  wire  s2_clock; // @[Cache.scala 476:18]
  wire  s2_reset; // @[Cache.scala 476:18]
  wire  s2_io_in_ready; // @[Cache.scala 476:18]
  wire  s2_io_in_valid; // @[Cache.scala 476:18]
  wire [31:0] s2_io_in_bits_req_addr; // @[Cache.scala 476:18]
  wire [2:0] s2_io_in_bits_req_size; // @[Cache.scala 476:18]
  wire [3:0] s2_io_in_bits_req_cmd; // @[Cache.scala 476:18]
  wire [7:0] s2_io_in_bits_req_wmask; // @[Cache.scala 476:18]
  wire [63:0] s2_io_in_bits_req_wdata; // @[Cache.scala 476:18]
  wire  s2_io_out_ready; // @[Cache.scala 476:18]
  wire  s2_io_out_valid; // @[Cache.scala 476:18]
  wire [31:0] s2_io_out_bits_req_addr; // @[Cache.scala 476:18]
  wire [2:0] s2_io_out_bits_req_size; // @[Cache.scala 476:18]
  wire [3:0] s2_io_out_bits_req_cmd; // @[Cache.scala 476:18]
  wire [7:0] s2_io_out_bits_req_wmask; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_req_wdata; // @[Cache.scala 476:18]
  wire [18:0] s2_io_out_bits_metas_0_tag; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_0_valid; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_0_dirty; // @[Cache.scala 476:18]
  wire [18:0] s2_io_out_bits_metas_1_tag; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_1_valid; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_1_dirty; // @[Cache.scala 476:18]
  wire [18:0] s2_io_out_bits_metas_2_tag; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_2_valid; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_2_dirty; // @[Cache.scala 476:18]
  wire [18:0] s2_io_out_bits_metas_3_tag; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_3_valid; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_3_dirty; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_datas_0_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_datas_1_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_datas_2_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_datas_3_data; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_hit; // @[Cache.scala 476:18]
  wire [3:0] s2_io_out_bits_waymask; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_mmio; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_isForwardData; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_forwardData_data_data; // @[Cache.scala 476:18]
  wire [3:0] s2_io_out_bits_forwardData_waymask; // @[Cache.scala 476:18]
  wire [18:0] s2_io_metaReadResp_0_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_0_valid; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_0_dirty; // @[Cache.scala 476:18]
  wire [18:0] s2_io_metaReadResp_1_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_1_valid; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_1_dirty; // @[Cache.scala 476:18]
  wire [18:0] s2_io_metaReadResp_2_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_2_valid; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_2_dirty; // @[Cache.scala 476:18]
  wire [18:0] s2_io_metaReadResp_3_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_3_valid; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_3_dirty; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataReadResp_0_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataReadResp_1_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataReadResp_2_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataReadResp_3_data; // @[Cache.scala 476:18]
  wire  s2_io_metaWriteBus_req_valid; // @[Cache.scala 476:18]
  wire [6:0] s2_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 476:18]
  wire [18:0] s2_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 476:18]
  wire [3:0] s2_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 476:18]
  wire  s2_io_dataWriteBus_req_valid; // @[Cache.scala 476:18]
  wire [9:0] s2_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 476:18]
  wire [3:0] s2_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 476:18]
  wire  s3_clock; // @[Cache.scala 477:18]
  wire  s3_reset; // @[Cache.scala 477:18]
  wire  s3_io_in_ready; // @[Cache.scala 477:18]
  wire  s3_io_in_valid; // @[Cache.scala 477:18]
  wire [31:0] s3_io_in_bits_req_addr; // @[Cache.scala 477:18]
  wire [2:0] s3_io_in_bits_req_size; // @[Cache.scala 477:18]
  wire [3:0] s3_io_in_bits_req_cmd; // @[Cache.scala 477:18]
  wire [7:0] s3_io_in_bits_req_wmask; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_req_wdata; // @[Cache.scala 477:18]
  wire [18:0] s3_io_in_bits_metas_0_tag; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_0_valid; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_0_dirty; // @[Cache.scala 477:18]
  wire [18:0] s3_io_in_bits_metas_1_tag; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_1_valid; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_1_dirty; // @[Cache.scala 477:18]
  wire [18:0] s3_io_in_bits_metas_2_tag; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_2_valid; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_2_dirty; // @[Cache.scala 477:18]
  wire [18:0] s3_io_in_bits_metas_3_tag; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_3_valid; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_3_dirty; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_datas_0_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_datas_1_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_datas_2_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_datas_3_data; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_hit; // @[Cache.scala 477:18]
  wire [3:0] s3_io_in_bits_waymask; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_mmio; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_isForwardData; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_forwardData_data_data; // @[Cache.scala 477:18]
  wire [3:0] s3_io_in_bits_forwardData_waymask; // @[Cache.scala 477:18]
  wire  s3_io_out_ready; // @[Cache.scala 477:18]
  wire  s3_io_out_valid; // @[Cache.scala 477:18]
  wire [3:0] s3_io_out_bits_cmd; // @[Cache.scala 477:18]
  wire [63:0] s3_io_out_bits_rdata; // @[Cache.scala 477:18]
  wire  s3_io_isFinish; // @[Cache.scala 477:18]
  wire  s3_io_dataReadBus_req_ready; // @[Cache.scala 477:18]
  wire  s3_io_dataReadBus_req_valid; // @[Cache.scala 477:18]
  wire [9:0] s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataReadBus_resp_data_0_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataReadBus_resp_data_1_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataReadBus_resp_data_2_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataReadBus_resp_data_3_data; // @[Cache.scala 477:18]
  wire  s3_io_dataWriteBus_req_valid; // @[Cache.scala 477:18]
  wire [9:0] s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 477:18]
  wire [3:0] s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 477:18]
  wire  s3_io_metaWriteBus_req_valid; // @[Cache.scala 477:18]
  wire [6:0] s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 477:18]
  wire [18:0] s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 477:18]
  wire  s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 477:18]
  wire [3:0] s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 477:18]
  wire  s3_io_mem_req_ready; // @[Cache.scala 477:18]
  wire  s3_io_mem_req_valid; // @[Cache.scala 477:18]
  wire [31:0] s3_io_mem_req_bits_addr; // @[Cache.scala 477:18]
  wire [3:0] s3_io_mem_req_bits_cmd; // @[Cache.scala 477:18]
  wire [63:0] s3_io_mem_req_bits_wdata; // @[Cache.scala 477:18]
  wire  s3_io_mem_resp_ready; // @[Cache.scala 477:18]
  wire  s3_io_mem_resp_valid; // @[Cache.scala 477:18]
  wire [3:0] s3_io_mem_resp_bits_cmd; // @[Cache.scala 477:18]
  wire [63:0] s3_io_mem_resp_bits_rdata; // @[Cache.scala 477:18]
  wire  s3_io_mmio_req_ready; // @[Cache.scala 477:18]
  wire  s3_io_mmio_req_valid; // @[Cache.scala 477:18]
  wire [31:0] s3_io_mmio_req_bits_addr; // @[Cache.scala 477:18]
  wire [2:0] s3_io_mmio_req_bits_size; // @[Cache.scala 477:18]
  wire [3:0] s3_io_mmio_req_bits_cmd; // @[Cache.scala 477:18]
  wire [7:0] s3_io_mmio_req_bits_wmask; // @[Cache.scala 477:18]
  wire [63:0] s3_io_mmio_req_bits_wdata; // @[Cache.scala 477:18]
  wire  s3_io_mmio_resp_ready; // @[Cache.scala 477:18]
  wire  s3_io_mmio_resp_valid; // @[Cache.scala 477:18]
  wire [63:0] s3_io_mmio_resp_bits_rdata; // @[Cache.scala 477:18]
  wire  s3_io_cohResp_valid; // @[Cache.scala 477:18]
  wire [3:0] s3_io_cohResp_bits_cmd; // @[Cache.scala 477:18]
  wire [63:0] s3_io_cohResp_bits_rdata; // @[Cache.scala 477:18]
  wire  s3_io_dataReadRespToL1; // @[Cache.scala 477:18]
  wire  metaArray_clock; // @[Cache.scala 478:25]
  wire  metaArray_reset; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_req_ready; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_req_valid; // @[Cache.scala 478:25]
  wire [6:0] metaArray_io_r0_req_bits_setIdx; // @[Cache.scala 478:25]
  wire [18:0] metaArray_io_r0_resp_data_0_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_resp_data_0_valid; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_resp_data_0_dirty; // @[Cache.scala 478:25]
  wire [18:0] metaArray_io_r0_resp_data_1_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_resp_data_1_valid; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_resp_data_1_dirty; // @[Cache.scala 478:25]
  wire [18:0] metaArray_io_r0_resp_data_2_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_resp_data_2_valid; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_resp_data_2_dirty; // @[Cache.scala 478:25]
  wire [18:0] metaArray_io_r0_resp_data_3_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_resp_data_3_valid; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_resp_data_3_dirty; // @[Cache.scala 478:25]
  wire  metaArray_io_wreq_valid; // @[Cache.scala 478:25]
  wire [6:0] metaArray_io_wreq_bits_setIdx; // @[Cache.scala 478:25]
  wire [18:0] metaArray_io_wreq_bits_data_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_wreq_bits_data_dirty; // @[Cache.scala 478:25]
  wire [3:0] metaArray_io_wreq_bits_waymask; // @[Cache.scala 478:25]
  wire  dataArray_clock; // @[Cache.scala 479:25]
  wire  dataArray_reset; // @[Cache.scala 479:25]
  wire  dataArray_io_r0_req_ready; // @[Cache.scala 479:25]
  wire  dataArray_io_r0_req_valid; // @[Cache.scala 479:25]
  wire [9:0] dataArray_io_r0_req_bits_setIdx; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r0_resp_data_0_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r0_resp_data_1_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r0_resp_data_2_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r0_resp_data_3_data; // @[Cache.scala 479:25]
  wire  dataArray_io_r1_req_ready; // @[Cache.scala 479:25]
  wire  dataArray_io_r1_req_valid; // @[Cache.scala 479:25]
  wire [9:0] dataArray_io_r1_req_bits_setIdx; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r1_resp_data_0_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r1_resp_data_1_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r1_resp_data_2_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r1_resp_data_3_data; // @[Cache.scala 479:25]
  wire  dataArray_io_wreq_valid; // @[Cache.scala 479:25]
  wire [9:0] dataArray_io_wreq_bits_setIdx; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_wreq_bits_data_data; // @[Cache.scala 479:25]
  wire [3:0] dataArray_io_wreq_bits_waymask; // @[Cache.scala 479:25]
  wire  arb_io_in_0_ready; // @[Cache.scala 488:19]
  wire  arb_io_in_0_valid; // @[Cache.scala 488:19]
  wire [31:0] arb_io_in_0_bits_addr; // @[Cache.scala 488:19]
  wire [2:0] arb_io_in_0_bits_size; // @[Cache.scala 488:19]
  wire [3:0] arb_io_in_0_bits_cmd; // @[Cache.scala 488:19]
  wire [7:0] arb_io_in_0_bits_wmask; // @[Cache.scala 488:19]
  wire [63:0] arb_io_in_0_bits_wdata; // @[Cache.scala 488:19]
  wire  arb_io_in_1_ready; // @[Cache.scala 488:19]
  wire  arb_io_in_1_valid; // @[Cache.scala 488:19]
  wire [31:0] arb_io_in_1_bits_addr; // @[Cache.scala 488:19]
  wire [2:0] arb_io_in_1_bits_size; // @[Cache.scala 488:19]
  wire [3:0] arb_io_in_1_bits_cmd; // @[Cache.scala 488:19]
  wire [7:0] arb_io_in_1_bits_wmask; // @[Cache.scala 488:19]
  wire [63:0] arb_io_in_1_bits_wdata; // @[Cache.scala 488:19]
  wire  arb_io_out_ready; // @[Cache.scala 488:19]
  wire  arb_io_out_valid; // @[Cache.scala 488:19]
  wire [31:0] arb_io_out_bits_addr; // @[Cache.scala 488:19]
  wire [2:0] arb_io_out_bits_size; // @[Cache.scala 488:19]
  wire [3:0] arb_io_out_bits_cmd; // @[Cache.scala 488:19]
  wire [7:0] arb_io_out_bits_wmask; // @[Cache.scala 488:19]
  wire [63:0] arb_io_out_bits_wdata; // @[Cache.scala 488:19]
  wire  _T = s2_io_out_ready & s2_io_out_valid; // @[Decoupled.scala 40:37]
  reg  _T_2; // @[Pipeline.scala 24:24]
  wire  _GEN_0 = _T ? 1'h0 : _T_2; // @[Pipeline.scala 25:25]
  wire  _T_3 = s1_io_out_valid & s2_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_1 = _T_3 | _GEN_0; // @[Pipeline.scala 26:38]
  reg [31:0] _T_5_req_addr; // @[Reg.scala 15:16]
  reg [2:0] _T_5_req_size; // @[Reg.scala 15:16]
  reg [3:0] _T_5_req_cmd; // @[Reg.scala 15:16]
  reg [7:0] _T_5_req_wmask; // @[Reg.scala 15:16]
  reg [63:0] _T_5_req_wdata; // @[Reg.scala 15:16]
  reg  _T_7; // @[Pipeline.scala 24:24]
  wire  _GEN_8 = s3_io_isFinish ? 1'h0 : _T_7; // @[Pipeline.scala 25:25]
  wire  _T_8 = s2_io_out_valid & s3_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_9 = _T_8 | _GEN_8; // @[Pipeline.scala 26:38]
  reg [31:0] _T_10_req_addr; // @[Reg.scala 15:16]
  reg [2:0] _T_10_req_size; // @[Reg.scala 15:16]
  reg [3:0] _T_10_req_cmd; // @[Reg.scala 15:16]
  reg [7:0] _T_10_req_wmask; // @[Reg.scala 15:16]
  reg [63:0] _T_10_req_wdata; // @[Reg.scala 15:16]
  reg [18:0] _T_10_metas_0_tag; // @[Reg.scala 15:16]
  reg  _T_10_metas_0_valid; // @[Reg.scala 15:16]
  reg  _T_10_metas_0_dirty; // @[Reg.scala 15:16]
  reg [18:0] _T_10_metas_1_tag; // @[Reg.scala 15:16]
  reg  _T_10_metas_1_valid; // @[Reg.scala 15:16]
  reg  _T_10_metas_1_dirty; // @[Reg.scala 15:16]
  reg [18:0] _T_10_metas_2_tag; // @[Reg.scala 15:16]
  reg  _T_10_metas_2_valid; // @[Reg.scala 15:16]
  reg  _T_10_metas_2_dirty; // @[Reg.scala 15:16]
  reg [18:0] _T_10_metas_3_tag; // @[Reg.scala 15:16]
  reg  _T_10_metas_3_valid; // @[Reg.scala 15:16]
  reg  _T_10_metas_3_dirty; // @[Reg.scala 15:16]
  reg [63:0] _T_10_datas_0_data; // @[Reg.scala 15:16]
  reg [63:0] _T_10_datas_1_data; // @[Reg.scala 15:16]
  reg [63:0] _T_10_datas_2_data; // @[Reg.scala 15:16]
  reg [63:0] _T_10_datas_3_data; // @[Reg.scala 15:16]
  reg  _T_10_hit; // @[Reg.scala 15:16]
  reg [3:0] _T_10_waymask; // @[Reg.scala 15:16]
  reg  _T_10_mmio; // @[Reg.scala 15:16]
  reg  _T_10_isForwardData; // @[Reg.scala 15:16]
  reg [63:0] _T_10_forwardData_data_data; // @[Reg.scala 15:16]
  reg [3:0] _T_10_forwardData_waymask; // @[Reg.scala 15:16]
  wire  _T_15 = s3_io_out_bits_cmd == 4'h4; // @[SimpleBus.scala 95:26]
  wire  _T_16 = s3_io_out_valid & _T_15; // @[Cache.scala 505:43]
  wire  _T_17 = s3_io_out_valid | s3_io_dataReadRespToL1; // @[Cache.scala 505:100]
  CacheStage1_1 s1 ( // @[Cache.scala 475:18]
    .io_in_ready(s1_io_in_ready),
    .io_in_valid(s1_io_in_valid),
    .io_in_bits_addr(s1_io_in_bits_addr),
    .io_in_bits_size(s1_io_in_bits_size),
    .io_in_bits_cmd(s1_io_in_bits_cmd),
    .io_in_bits_wmask(s1_io_in_bits_wmask),
    .io_in_bits_wdata(s1_io_in_bits_wdata),
    .io_out_ready(s1_io_out_ready),
    .io_out_valid(s1_io_out_valid),
    .io_out_bits_req_addr(s1_io_out_bits_req_addr),
    .io_out_bits_req_size(s1_io_out_bits_req_size),
    .io_out_bits_req_cmd(s1_io_out_bits_req_cmd),
    .io_out_bits_req_wmask(s1_io_out_bits_req_wmask),
    .io_out_bits_req_wdata(s1_io_out_bits_req_wdata),
    .io_metaReadBus_req_ready(s1_io_metaReadBus_req_ready),
    .io_metaReadBus_req_valid(s1_io_metaReadBus_req_valid),
    .io_metaReadBus_req_bits_setIdx(s1_io_metaReadBus_req_bits_setIdx),
    .io_metaReadBus_resp_data_0_tag(s1_io_metaReadBus_resp_data_0_tag),
    .io_metaReadBus_resp_data_0_valid(s1_io_metaReadBus_resp_data_0_valid),
    .io_metaReadBus_resp_data_0_dirty(s1_io_metaReadBus_resp_data_0_dirty),
    .io_metaReadBus_resp_data_1_tag(s1_io_metaReadBus_resp_data_1_tag),
    .io_metaReadBus_resp_data_1_valid(s1_io_metaReadBus_resp_data_1_valid),
    .io_metaReadBus_resp_data_1_dirty(s1_io_metaReadBus_resp_data_1_dirty),
    .io_metaReadBus_resp_data_2_tag(s1_io_metaReadBus_resp_data_2_tag),
    .io_metaReadBus_resp_data_2_valid(s1_io_metaReadBus_resp_data_2_valid),
    .io_metaReadBus_resp_data_2_dirty(s1_io_metaReadBus_resp_data_2_dirty),
    .io_metaReadBus_resp_data_3_tag(s1_io_metaReadBus_resp_data_3_tag),
    .io_metaReadBus_resp_data_3_valid(s1_io_metaReadBus_resp_data_3_valid),
    .io_metaReadBus_resp_data_3_dirty(s1_io_metaReadBus_resp_data_3_dirty),
    .io_dataReadBus_req_ready(s1_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s1_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s1_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s1_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s1_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s1_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s1_io_dataReadBus_resp_data_3_data)
  );
  CacheStage2_1 s2 ( // @[Cache.scala 476:18]
    .clock(s2_clock),
    .reset(s2_reset),
    .io_in_ready(s2_io_in_ready),
    .io_in_valid(s2_io_in_valid),
    .io_in_bits_req_addr(s2_io_in_bits_req_addr),
    .io_in_bits_req_size(s2_io_in_bits_req_size),
    .io_in_bits_req_cmd(s2_io_in_bits_req_cmd),
    .io_in_bits_req_wmask(s2_io_in_bits_req_wmask),
    .io_in_bits_req_wdata(s2_io_in_bits_req_wdata),
    .io_out_ready(s2_io_out_ready),
    .io_out_valid(s2_io_out_valid),
    .io_out_bits_req_addr(s2_io_out_bits_req_addr),
    .io_out_bits_req_size(s2_io_out_bits_req_size),
    .io_out_bits_req_cmd(s2_io_out_bits_req_cmd),
    .io_out_bits_req_wmask(s2_io_out_bits_req_wmask),
    .io_out_bits_req_wdata(s2_io_out_bits_req_wdata),
    .io_out_bits_metas_0_tag(s2_io_out_bits_metas_0_tag),
    .io_out_bits_metas_0_valid(s2_io_out_bits_metas_0_valid),
    .io_out_bits_metas_0_dirty(s2_io_out_bits_metas_0_dirty),
    .io_out_bits_metas_1_tag(s2_io_out_bits_metas_1_tag),
    .io_out_bits_metas_1_valid(s2_io_out_bits_metas_1_valid),
    .io_out_bits_metas_1_dirty(s2_io_out_bits_metas_1_dirty),
    .io_out_bits_metas_2_tag(s2_io_out_bits_metas_2_tag),
    .io_out_bits_metas_2_valid(s2_io_out_bits_metas_2_valid),
    .io_out_bits_metas_2_dirty(s2_io_out_bits_metas_2_dirty),
    .io_out_bits_metas_3_tag(s2_io_out_bits_metas_3_tag),
    .io_out_bits_metas_3_valid(s2_io_out_bits_metas_3_valid),
    .io_out_bits_metas_3_dirty(s2_io_out_bits_metas_3_dirty),
    .io_out_bits_datas_0_data(s2_io_out_bits_datas_0_data),
    .io_out_bits_datas_1_data(s2_io_out_bits_datas_1_data),
    .io_out_bits_datas_2_data(s2_io_out_bits_datas_2_data),
    .io_out_bits_datas_3_data(s2_io_out_bits_datas_3_data),
    .io_out_bits_hit(s2_io_out_bits_hit),
    .io_out_bits_waymask(s2_io_out_bits_waymask),
    .io_out_bits_mmio(s2_io_out_bits_mmio),
    .io_out_bits_isForwardData(s2_io_out_bits_isForwardData),
    .io_out_bits_forwardData_data_data(s2_io_out_bits_forwardData_data_data),
    .io_out_bits_forwardData_waymask(s2_io_out_bits_forwardData_waymask),
    .io_metaReadResp_0_tag(s2_io_metaReadResp_0_tag),
    .io_metaReadResp_0_valid(s2_io_metaReadResp_0_valid),
    .io_metaReadResp_0_dirty(s2_io_metaReadResp_0_dirty),
    .io_metaReadResp_1_tag(s2_io_metaReadResp_1_tag),
    .io_metaReadResp_1_valid(s2_io_metaReadResp_1_valid),
    .io_metaReadResp_1_dirty(s2_io_metaReadResp_1_dirty),
    .io_metaReadResp_2_tag(s2_io_metaReadResp_2_tag),
    .io_metaReadResp_2_valid(s2_io_metaReadResp_2_valid),
    .io_metaReadResp_2_dirty(s2_io_metaReadResp_2_dirty),
    .io_metaReadResp_3_tag(s2_io_metaReadResp_3_tag),
    .io_metaReadResp_3_valid(s2_io_metaReadResp_3_valid),
    .io_metaReadResp_3_dirty(s2_io_metaReadResp_3_dirty),
    .io_dataReadResp_0_data(s2_io_dataReadResp_0_data),
    .io_dataReadResp_1_data(s2_io_dataReadResp_1_data),
    .io_dataReadResp_2_data(s2_io_dataReadResp_2_data),
    .io_dataReadResp_3_data(s2_io_dataReadResp_3_data),
    .io_metaWriteBus_req_valid(s2_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s2_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s2_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_dirty(s2_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s2_io_metaWriteBus_req_bits_waymask),
    .io_dataWriteBus_req_valid(s2_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s2_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s2_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s2_io_dataWriteBus_req_bits_waymask)
  );
  CacheStage3_1 s3 ( // @[Cache.scala 477:18]
    .clock(s3_clock),
    .reset(s3_reset),
    .io_in_ready(s3_io_in_ready),
    .io_in_valid(s3_io_in_valid),
    .io_in_bits_req_addr(s3_io_in_bits_req_addr),
    .io_in_bits_req_size(s3_io_in_bits_req_size),
    .io_in_bits_req_cmd(s3_io_in_bits_req_cmd),
    .io_in_bits_req_wmask(s3_io_in_bits_req_wmask),
    .io_in_bits_req_wdata(s3_io_in_bits_req_wdata),
    .io_in_bits_metas_0_tag(s3_io_in_bits_metas_0_tag),
    .io_in_bits_metas_0_valid(s3_io_in_bits_metas_0_valid),
    .io_in_bits_metas_0_dirty(s3_io_in_bits_metas_0_dirty),
    .io_in_bits_metas_1_tag(s3_io_in_bits_metas_1_tag),
    .io_in_bits_metas_1_valid(s3_io_in_bits_metas_1_valid),
    .io_in_bits_metas_1_dirty(s3_io_in_bits_metas_1_dirty),
    .io_in_bits_metas_2_tag(s3_io_in_bits_metas_2_tag),
    .io_in_bits_metas_2_valid(s3_io_in_bits_metas_2_valid),
    .io_in_bits_metas_2_dirty(s3_io_in_bits_metas_2_dirty),
    .io_in_bits_metas_3_tag(s3_io_in_bits_metas_3_tag),
    .io_in_bits_metas_3_valid(s3_io_in_bits_metas_3_valid),
    .io_in_bits_metas_3_dirty(s3_io_in_bits_metas_3_dirty),
    .io_in_bits_datas_0_data(s3_io_in_bits_datas_0_data),
    .io_in_bits_datas_1_data(s3_io_in_bits_datas_1_data),
    .io_in_bits_datas_2_data(s3_io_in_bits_datas_2_data),
    .io_in_bits_datas_3_data(s3_io_in_bits_datas_3_data),
    .io_in_bits_hit(s3_io_in_bits_hit),
    .io_in_bits_waymask(s3_io_in_bits_waymask),
    .io_in_bits_mmio(s3_io_in_bits_mmio),
    .io_in_bits_isForwardData(s3_io_in_bits_isForwardData),
    .io_in_bits_forwardData_data_data(s3_io_in_bits_forwardData_data_data),
    .io_in_bits_forwardData_waymask(s3_io_in_bits_forwardData_waymask),
    .io_out_ready(s3_io_out_ready),
    .io_out_valid(s3_io_out_valid),
    .io_out_bits_cmd(s3_io_out_bits_cmd),
    .io_out_bits_rdata(s3_io_out_bits_rdata),
    .io_isFinish(s3_io_isFinish),
    .io_dataReadBus_req_ready(s3_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s3_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s3_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s3_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s3_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s3_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s3_io_dataReadBus_resp_data_3_data),
    .io_dataWriteBus_req_valid(s3_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s3_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s3_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s3_io_dataWriteBus_req_bits_waymask),
    .io_metaWriteBus_req_valid(s3_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s3_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s3_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_dirty(s3_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s3_io_metaWriteBus_req_bits_waymask),
    .io_mem_req_ready(s3_io_mem_req_ready),
    .io_mem_req_valid(s3_io_mem_req_valid),
    .io_mem_req_bits_addr(s3_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(s3_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(s3_io_mem_req_bits_wdata),
    .io_mem_resp_ready(s3_io_mem_resp_ready),
    .io_mem_resp_valid(s3_io_mem_resp_valid),
    .io_mem_resp_bits_cmd(s3_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_rdata(s3_io_mem_resp_bits_rdata),
    .io_mmio_req_ready(s3_io_mmio_req_ready),
    .io_mmio_req_valid(s3_io_mmio_req_valid),
    .io_mmio_req_bits_addr(s3_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size(s3_io_mmio_req_bits_size),
    .io_mmio_req_bits_cmd(s3_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(s3_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(s3_io_mmio_req_bits_wdata),
    .io_mmio_resp_ready(s3_io_mmio_resp_ready),
    .io_mmio_resp_valid(s3_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(s3_io_mmio_resp_bits_rdata),
    .io_cohResp_valid(s3_io_cohResp_valid),
    .io_cohResp_bits_cmd(s3_io_cohResp_bits_cmd),
    .io_cohResp_bits_rdata(s3_io_cohResp_bits_rdata),
    .io_dataReadRespToL1(s3_io_dataReadRespToL1)
  );
  SRAMTemplateWithArbiter metaArray ( // @[Cache.scala 478:25]
    .clock(metaArray_clock),
    .reset(metaArray_reset),
    .io_r0_req_ready(metaArray_io_r0_req_ready),
    .io_r0_req_valid(metaArray_io_r0_req_valid),
    .io_r0_req_bits_setIdx(metaArray_io_r0_req_bits_setIdx),
    .io_r0_resp_data_0_tag(metaArray_io_r0_resp_data_0_tag),
    .io_r0_resp_data_0_valid(metaArray_io_r0_resp_data_0_valid),
    .io_r0_resp_data_0_dirty(metaArray_io_r0_resp_data_0_dirty),
    .io_r0_resp_data_1_tag(metaArray_io_r0_resp_data_1_tag),
    .io_r0_resp_data_1_valid(metaArray_io_r0_resp_data_1_valid),
    .io_r0_resp_data_1_dirty(metaArray_io_r0_resp_data_1_dirty),
    .io_r0_resp_data_2_tag(metaArray_io_r0_resp_data_2_tag),
    .io_r0_resp_data_2_valid(metaArray_io_r0_resp_data_2_valid),
    .io_r0_resp_data_2_dirty(metaArray_io_r0_resp_data_2_dirty),
    .io_r0_resp_data_3_tag(metaArray_io_r0_resp_data_3_tag),
    .io_r0_resp_data_3_valid(metaArray_io_r0_resp_data_3_valid),
    .io_r0_resp_data_3_dirty(metaArray_io_r0_resp_data_3_dirty),
    .io_wreq_valid(metaArray_io_wreq_valid),
    .io_wreq_bits_setIdx(metaArray_io_wreq_bits_setIdx),
    .io_wreq_bits_data_tag(metaArray_io_wreq_bits_data_tag),
    .io_wreq_bits_data_dirty(metaArray_io_wreq_bits_data_dirty),
    .io_wreq_bits_waymask(metaArray_io_wreq_bits_waymask)
  );
  SRAMTemplateWithArbiter_1 dataArray ( // @[Cache.scala 479:25]
    .clock(dataArray_clock),
    .reset(dataArray_reset),
    .io_r0_req_ready(dataArray_io_r0_req_ready),
    .io_r0_req_valid(dataArray_io_r0_req_valid),
    .io_r0_req_bits_setIdx(dataArray_io_r0_req_bits_setIdx),
    .io_r0_resp_data_0_data(dataArray_io_r0_resp_data_0_data),
    .io_r0_resp_data_1_data(dataArray_io_r0_resp_data_1_data),
    .io_r0_resp_data_2_data(dataArray_io_r0_resp_data_2_data),
    .io_r0_resp_data_3_data(dataArray_io_r0_resp_data_3_data),
    .io_r1_req_ready(dataArray_io_r1_req_ready),
    .io_r1_req_valid(dataArray_io_r1_req_valid),
    .io_r1_req_bits_setIdx(dataArray_io_r1_req_bits_setIdx),
    .io_r1_resp_data_0_data(dataArray_io_r1_resp_data_0_data),
    .io_r1_resp_data_1_data(dataArray_io_r1_resp_data_1_data),
    .io_r1_resp_data_2_data(dataArray_io_r1_resp_data_2_data),
    .io_r1_resp_data_3_data(dataArray_io_r1_resp_data_3_data),
    .io_wreq_valid(dataArray_io_wreq_valid),
    .io_wreq_bits_setIdx(dataArray_io_wreq_bits_setIdx),
    .io_wreq_bits_data_data(dataArray_io_wreq_bits_data_data),
    .io_wreq_bits_waymask(dataArray_io_wreq_bits_waymask)
  );
  Arbiter_9 arb ( // @[Cache.scala 488:19]
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_addr(arb_io_in_0_bits_addr),
    .io_in_0_bits_size(arb_io_in_0_bits_size),
    .io_in_0_bits_cmd(arb_io_in_0_bits_cmd),
    .io_in_0_bits_wmask(arb_io_in_0_bits_wmask),
    .io_in_0_bits_wdata(arb_io_in_0_bits_wdata),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_addr(arb_io_in_1_bits_addr),
    .io_in_1_bits_size(arb_io_in_1_bits_size),
    .io_in_1_bits_cmd(arb_io_in_1_bits_cmd),
    .io_in_1_bits_wmask(arb_io_in_1_bits_wmask),
    .io_in_1_bits_wdata(arb_io_in_1_bits_wdata),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_addr(arb_io_out_bits_addr),
    .io_out_bits_size(arb_io_out_bits_size),
    .io_out_bits_cmd(arb_io_out_bits_cmd),
    .io_out_bits_wmask(arb_io_out_bits_wmask),
    .io_out_bits_wdata(arb_io_out_bits_wdata)
  );
  assign io_in_req_ready = arb_io_in_1_ready; // @[Cache.scala 489:28]
  assign io_in_resp_valid = _T_16 ? 1'h0 : _T_17; // @[Cache.scala 499:14 Cache.scala 505:20]
  assign io_in_resp_bits_cmd = s3_io_out_bits_cmd; // @[Cache.scala 499:14]
  assign io_in_resp_bits_rdata = s3_io_out_bits_rdata; // @[Cache.scala 499:14]
  assign io_out_mem_req_valid = s3_io_mem_req_valid; // @[Cache.scala 501:14]
  assign io_out_mem_req_bits_addr = s3_io_mem_req_bits_addr; // @[Cache.scala 501:14]
  assign io_out_mem_req_bits_cmd = s3_io_mem_req_bits_cmd; // @[Cache.scala 501:14]
  assign io_out_mem_req_bits_wdata = s3_io_mem_req_bits_wdata; // @[Cache.scala 501:14]
  assign io_out_coh_req_ready = arb_io_in_0_ready; // @[Cache.scala 514:26]
  assign io_out_coh_resp_valid = s3_io_cohResp_valid; // @[Cache.scala 515:21]
  assign io_out_coh_resp_bits_cmd = s3_io_cohResp_bits_cmd; // @[Cache.scala 515:21]
  assign io_out_coh_resp_bits_rdata = s3_io_cohResp_bits_rdata; // @[Cache.scala 515:21]
  assign io_mmio_req_valid = s3_io_mmio_req_valid; // @[Cache.scala 502:11]
  assign io_mmio_req_bits_addr = s3_io_mmio_req_bits_addr; // @[Cache.scala 502:11]
  assign io_mmio_req_bits_size = s3_io_mmio_req_bits_size; // @[Cache.scala 502:11]
  assign io_mmio_req_bits_cmd = s3_io_mmio_req_bits_cmd; // @[Cache.scala 502:11]
  assign io_mmio_req_bits_wmask = s3_io_mmio_req_bits_wmask; // @[Cache.scala 502:11]
  assign io_mmio_req_bits_wdata = s3_io_mmio_req_bits_wdata; // @[Cache.scala 502:11]
  assign s1_io_in_valid = arb_io_out_valid; // @[Cache.scala 491:12]
  assign s1_io_in_bits_addr = arb_io_out_bits_addr; // @[Cache.scala 491:12]
  assign s1_io_in_bits_size = arb_io_out_bits_size; // @[Cache.scala 491:12]
  assign s1_io_in_bits_cmd = arb_io_out_bits_cmd; // @[Cache.scala 491:12]
  assign s1_io_in_bits_wmask = arb_io_out_bits_wmask; // @[Cache.scala 491:12]
  assign s1_io_in_bits_wdata = arb_io_out_bits_wdata; // @[Cache.scala 491:12]
  assign s1_io_out_ready = s2_io_in_ready; // @[Pipeline.scala 29:16]
  assign s1_io_metaReadBus_req_ready = metaArray_io_r0_req_ready; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_0_tag = metaArray_io_r0_resp_data_0_tag; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_0_valid = metaArray_io_r0_resp_data_0_valid; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_0_dirty = metaArray_io_r0_resp_data_0_dirty; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_1_tag = metaArray_io_r0_resp_data_1_tag; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_1_valid = metaArray_io_r0_resp_data_1_valid; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_1_dirty = metaArray_io_r0_resp_data_1_dirty; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_2_tag = metaArray_io_r0_resp_data_2_tag; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_2_valid = metaArray_io_r0_resp_data_2_valid; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_2_dirty = metaArray_io_r0_resp_data_2_dirty; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_3_tag = metaArray_io_r0_resp_data_3_tag; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_3_valid = metaArray_io_r0_resp_data_3_valid; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_3_dirty = metaArray_io_r0_resp_data_3_dirty; // @[Cache.scala 523:21]
  assign s1_io_dataReadBus_req_ready = dataArray_io_r0_req_ready; // @[Cache.scala 524:21]
  assign s1_io_dataReadBus_resp_data_0_data = dataArray_io_r0_resp_data_0_data; // @[Cache.scala 524:21]
  assign s1_io_dataReadBus_resp_data_1_data = dataArray_io_r0_resp_data_1_data; // @[Cache.scala 524:21]
  assign s1_io_dataReadBus_resp_data_2_data = dataArray_io_r0_resp_data_2_data; // @[Cache.scala 524:21]
  assign s1_io_dataReadBus_resp_data_3_data = dataArray_io_r0_resp_data_3_data; // @[Cache.scala 524:21]
  assign s2_clock = clock;
  assign s2_reset = reset;
  assign s2_io_in_valid = _T_2; // @[Pipeline.scala 31:17]
  assign s2_io_in_bits_req_addr = _T_5_req_addr; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_size = _T_5_req_size; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_cmd = _T_5_req_cmd; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_wmask = _T_5_req_wmask; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_wdata = _T_5_req_wdata; // @[Pipeline.scala 30:16]
  assign s2_io_out_ready = s3_io_in_ready; // @[Pipeline.scala 29:16]
  assign s2_io_metaReadResp_0_tag = s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_0_valid = s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_0_dirty = s1_io_metaReadBus_resp_data_0_dirty; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_1_tag = s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_1_valid = s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_1_dirty = s1_io_metaReadBus_resp_data_1_dirty; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_2_tag = s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_2_valid = s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_2_dirty = s1_io_metaReadBus_resp_data_2_dirty; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_3_tag = s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_3_valid = s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_3_dirty = s1_io_metaReadBus_resp_data_3_dirty; // @[Cache.scala 530:22]
  assign s2_io_dataReadResp_0_data = s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 531:22]
  assign s2_io_dataReadResp_1_data = s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 531:22]
  assign s2_io_dataReadResp_2_data = s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 531:22]
  assign s2_io_dataReadResp_3_data = s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 531:22]
  assign s2_io_metaWriteBus_req_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 533:22]
  assign s2_io_metaWriteBus_req_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 533:22]
  assign s2_io_metaWriteBus_req_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 533:22]
  assign s2_io_metaWriteBus_req_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 533:22]
  assign s2_io_metaWriteBus_req_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 533:22]
  assign s2_io_dataWriteBus_req_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 532:22]
  assign s2_io_dataWriteBus_req_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 532:22]
  assign s2_io_dataWriteBus_req_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 532:22]
  assign s2_io_dataWriteBus_req_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 532:22]
  assign s3_clock = clock;
  assign s3_reset = reset;
  assign s3_io_in_valid = _T_7; // @[Pipeline.scala 31:17]
  assign s3_io_in_bits_req_addr = _T_10_req_addr; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_size = _T_10_req_size; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_cmd = _T_10_req_cmd; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_wmask = _T_10_req_wmask; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_wdata = _T_10_req_wdata; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_tag = _T_10_metas_0_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_valid = _T_10_metas_0_valid; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_dirty = _T_10_metas_0_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_tag = _T_10_metas_1_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_valid = _T_10_metas_1_valid; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_dirty = _T_10_metas_1_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_tag = _T_10_metas_2_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_valid = _T_10_metas_2_valid; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_dirty = _T_10_metas_2_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_tag = _T_10_metas_3_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_valid = _T_10_metas_3_valid; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_dirty = _T_10_metas_3_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_0_data = _T_10_datas_0_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_1_data = _T_10_datas_1_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_2_data = _T_10_datas_2_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_3_data = _T_10_datas_3_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_hit = _T_10_hit; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_waymask = _T_10_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_mmio = _T_10_mmio; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_isForwardData = _T_10_isForwardData; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_data_data = _T_10_forwardData_data_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_waymask = _T_10_forwardData_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_out_ready = io_in_resp_ready; // @[Cache.scala 499:14]
  assign s3_io_dataReadBus_req_ready = dataArray_io_r1_req_ready; // @[Cache.scala 525:21]
  assign s3_io_dataReadBus_resp_data_0_data = dataArray_io_r1_resp_data_0_data; // @[Cache.scala 525:21]
  assign s3_io_dataReadBus_resp_data_1_data = dataArray_io_r1_resp_data_1_data; // @[Cache.scala 525:21]
  assign s3_io_dataReadBus_resp_data_2_data = dataArray_io_r1_resp_data_2_data; // @[Cache.scala 525:21]
  assign s3_io_dataReadBus_resp_data_3_data = dataArray_io_r1_resp_data_3_data; // @[Cache.scala 525:21]
  assign s3_io_mem_req_ready = io_out_mem_req_ready; // @[Cache.scala 501:14]
  assign s3_io_mem_resp_valid = io_out_mem_resp_valid; // @[Cache.scala 501:14]
  assign s3_io_mem_resp_bits_cmd = io_out_mem_resp_bits_cmd; // @[Cache.scala 501:14]
  assign s3_io_mem_resp_bits_rdata = io_out_mem_resp_bits_rdata; // @[Cache.scala 501:14]
  assign s3_io_mmio_req_ready = io_mmio_req_ready; // @[Cache.scala 502:11]
  assign s3_io_mmio_resp_valid = io_mmio_resp_valid; // @[Cache.scala 502:11]
  assign s3_io_mmio_resp_bits_rdata = io_mmio_resp_bits_rdata; // @[Cache.scala 502:11]
  assign metaArray_clock = clock;
  assign metaArray_reset = reset;
  assign metaArray_io_r0_req_valid = s1_io_metaReadBus_req_valid; // @[Cache.scala 523:21]
  assign metaArray_io_r0_req_bits_setIdx = s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 523:21]
  assign metaArray_io_wreq_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 527:18]
  assign metaArray_io_wreq_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 527:18]
  assign metaArray_io_wreq_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 527:18]
  assign metaArray_io_wreq_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 527:18]
  assign metaArray_io_wreq_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 527:18]
  assign dataArray_clock = clock;
  assign dataArray_reset = reset;
  assign dataArray_io_r0_req_valid = s1_io_dataReadBus_req_valid; // @[Cache.scala 524:21]
  assign dataArray_io_r0_req_bits_setIdx = s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 524:21]
  assign dataArray_io_r1_req_valid = s3_io_dataReadBus_req_valid; // @[Cache.scala 525:21]
  assign dataArray_io_r1_req_bits_setIdx = s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 525:21]
  assign dataArray_io_wreq_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 528:18]
  assign dataArray_io_wreq_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 528:18]
  assign dataArray_io_wreq_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 528:18]
  assign dataArray_io_wreq_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 528:18]
  assign arb_io_in_0_valid = io_out_coh_req_valid; // @[Cache.scala 513:24]
  assign arb_io_in_0_bits_addr = io_out_coh_req_bits_addr; // @[Cache.scala 512:23]
  assign arb_io_in_0_bits_size = 3'h3; // @[Cache.scala 512:23]
  assign arb_io_in_0_bits_cmd = 4'h8; // @[Cache.scala 512:23]
  assign arb_io_in_0_bits_wmask = 8'hff; // @[Cache.scala 512:23]
  assign arb_io_in_0_bits_wdata = io_out_coh_req_bits_wdata; // @[Cache.scala 512:23]
  assign arb_io_in_1_valid = io_in_req_valid; // @[Cache.scala 489:28]
  assign arb_io_in_1_bits_addr = io_in_req_bits_addr; // @[Cache.scala 489:28]
  assign arb_io_in_1_bits_size = io_in_req_bits_size; // @[Cache.scala 489:28]
  assign arb_io_in_1_bits_cmd = io_in_req_bits_cmd; // @[Cache.scala 489:28]
  assign arb_io_in_1_bits_wmask = io_in_req_bits_wmask; // @[Cache.scala 489:28]
  assign arb_io_in_1_bits_wdata = io_in_req_bits_wdata; // @[Cache.scala 489:28]
  assign arb_io_out_ready = s1_io_in_ready; // @[Cache.scala 491:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _T_5_req_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_5_req_size = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  _T_5_req_cmd = _RAND_3[3:0];
  _RAND_4 = {1{`RANDOM}};
  _T_5_req_wmask = _RAND_4[7:0];
  _RAND_5 = {2{`RANDOM}};
  _T_5_req_wdata = _RAND_5[63:0];
  _RAND_6 = {1{`RANDOM}};
  _T_7 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_10_req_addr = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  _T_10_req_size = _RAND_8[2:0];
  _RAND_9 = {1{`RANDOM}};
  _T_10_req_cmd = _RAND_9[3:0];
  _RAND_10 = {1{`RANDOM}};
  _T_10_req_wmask = _RAND_10[7:0];
  _RAND_11 = {2{`RANDOM}};
  _T_10_req_wdata = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  _T_10_metas_0_tag = _RAND_12[18:0];
  _RAND_13 = {1{`RANDOM}};
  _T_10_metas_0_valid = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _T_10_metas_0_dirty = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _T_10_metas_1_tag = _RAND_15[18:0];
  _RAND_16 = {1{`RANDOM}};
  _T_10_metas_1_valid = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  _T_10_metas_1_dirty = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _T_10_metas_2_tag = _RAND_18[18:0];
  _RAND_19 = {1{`RANDOM}};
  _T_10_metas_2_valid = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  _T_10_metas_2_dirty = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _T_10_metas_3_tag = _RAND_21[18:0];
  _RAND_22 = {1{`RANDOM}};
  _T_10_metas_3_valid = _RAND_22[0:0];
  _RAND_23 = {1{`RANDOM}};
  _T_10_metas_3_dirty = _RAND_23[0:0];
  _RAND_24 = {2{`RANDOM}};
  _T_10_datas_0_data = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  _T_10_datas_1_data = _RAND_25[63:0];
  _RAND_26 = {2{`RANDOM}};
  _T_10_datas_2_data = _RAND_26[63:0];
  _RAND_27 = {2{`RANDOM}};
  _T_10_datas_3_data = _RAND_27[63:0];
  _RAND_28 = {1{`RANDOM}};
  _T_10_hit = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  _T_10_waymask = _RAND_29[3:0];
  _RAND_30 = {1{`RANDOM}};
  _T_10_mmio = _RAND_30[0:0];
  _RAND_31 = {1{`RANDOM}};
  _T_10_isForwardData = _RAND_31[0:0];
  _RAND_32 = {2{`RANDOM}};
  _T_10_forwardData_data_data = _RAND_32[63:0];
  _RAND_33 = {1{`RANDOM}};
  _T_10_forwardData_waymask = _RAND_33[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_2 <= 1'h0;
    end else begin
      _T_2 <= _GEN_1;
    end
    if (_T_3) begin
      _T_5_req_addr <= s1_io_out_bits_req_addr;
    end
    if (_T_3) begin
      _T_5_req_size <= s1_io_out_bits_req_size;
    end
    if (_T_3) begin
      _T_5_req_cmd <= s1_io_out_bits_req_cmd;
    end
    if (_T_3) begin
      _T_5_req_wmask <= s1_io_out_bits_req_wmask;
    end
    if (_T_3) begin
      _T_5_req_wdata <= s1_io_out_bits_req_wdata;
    end
    if (reset) begin
      _T_7 <= 1'h0;
    end else begin
      _T_7 <= _GEN_9;
    end
    if (_T_8) begin
      _T_10_req_addr <= s2_io_out_bits_req_addr;
    end
    if (_T_8) begin
      _T_10_req_size <= s2_io_out_bits_req_size;
    end
    if (_T_8) begin
      _T_10_req_cmd <= s2_io_out_bits_req_cmd;
    end
    if (_T_8) begin
      _T_10_req_wmask <= s2_io_out_bits_req_wmask;
    end
    if (_T_8) begin
      _T_10_req_wdata <= s2_io_out_bits_req_wdata;
    end
    if (_T_8) begin
      _T_10_metas_0_tag <= s2_io_out_bits_metas_0_tag;
    end
    if (_T_8) begin
      _T_10_metas_0_valid <= s2_io_out_bits_metas_0_valid;
    end
    if (_T_8) begin
      _T_10_metas_0_dirty <= s2_io_out_bits_metas_0_dirty;
    end
    if (_T_8) begin
      _T_10_metas_1_tag <= s2_io_out_bits_metas_1_tag;
    end
    if (_T_8) begin
      _T_10_metas_1_valid <= s2_io_out_bits_metas_1_valid;
    end
    if (_T_8) begin
      _T_10_metas_1_dirty <= s2_io_out_bits_metas_1_dirty;
    end
    if (_T_8) begin
      _T_10_metas_2_tag <= s2_io_out_bits_metas_2_tag;
    end
    if (_T_8) begin
      _T_10_metas_2_valid <= s2_io_out_bits_metas_2_valid;
    end
    if (_T_8) begin
      _T_10_metas_2_dirty <= s2_io_out_bits_metas_2_dirty;
    end
    if (_T_8) begin
      _T_10_metas_3_tag <= s2_io_out_bits_metas_3_tag;
    end
    if (_T_8) begin
      _T_10_metas_3_valid <= s2_io_out_bits_metas_3_valid;
    end
    if (_T_8) begin
      _T_10_metas_3_dirty <= s2_io_out_bits_metas_3_dirty;
    end
    if (_T_8) begin
      _T_10_datas_0_data <= s2_io_out_bits_datas_0_data;
    end
    if (_T_8) begin
      _T_10_datas_1_data <= s2_io_out_bits_datas_1_data;
    end
    if (_T_8) begin
      _T_10_datas_2_data <= s2_io_out_bits_datas_2_data;
    end
    if (_T_8) begin
      _T_10_datas_3_data <= s2_io_out_bits_datas_3_data;
    end
    if (_T_8) begin
      _T_10_hit <= s2_io_out_bits_hit;
    end
    if (_T_8) begin
      _T_10_waymask <= s2_io_out_bits_waymask;
    end
    if (_T_8) begin
      _T_10_mmio <= s2_io_out_bits_mmio;
    end
    if (_T_8) begin
      _T_10_isForwardData <= s2_io_out_bits_isForwardData;
    end
    if (_T_8) begin
      _T_10_forwardData_data_data <= s2_io_out_bits_forwardData_data_data;
    end
    if (_T_8) begin
      _T_10_forwardData_waymask <= s2_io_out_bits_forwardData_waymask;
    end
  end
endmodule
module NutCore(
  input         clock,
  input         reset,
  input         io_imem_mem_req_ready,
  output        io_imem_mem_req_valid,
  output [31:0] io_imem_mem_req_bits_addr,
  output [3:0]  io_imem_mem_req_bits_cmd,
  output [63:0] io_imem_mem_req_bits_wdata,
  input         io_imem_mem_resp_valid,
  input  [3:0]  io_imem_mem_resp_bits_cmd,
  input  [63:0] io_imem_mem_resp_bits_rdata,
  input         io_dmem_mem_req_ready,
  output        io_dmem_mem_req_valid,
  output [31:0] io_dmem_mem_req_bits_addr,
  output [3:0]  io_dmem_mem_req_bits_cmd,
  output [63:0] io_dmem_mem_req_bits_wdata,
  input         io_dmem_mem_resp_valid,
  input  [3:0]  io_dmem_mem_resp_bits_cmd,
  input  [63:0] io_dmem_mem_resp_bits_rdata,
  output        io_dmem_coh_req_ready,
  input         io_dmem_coh_req_valid,
  input  [31:0] io_dmem_coh_req_bits_addr,
  input  [63:0] io_dmem_coh_req_bits_wdata,
  output        io_dmem_coh_resp_valid,
  output [3:0]  io_dmem_coh_resp_bits_cmd,
  output [63:0] io_dmem_coh_resp_bits_rdata,
  input         io_mmio_req_ready,
  output        io_mmio_req_valid,
  output [31:0] io_mmio_req_bits_addr,
  output [2:0]  io_mmio_req_bits_size,
  output [3:0]  io_mmio_req_bits_cmd,
  output [7:0]  io_mmio_req_bits_wmask,
  output [63:0] io_mmio_req_bits_wdata,
  input         io_mmio_resp_valid,
  input  [3:0]  io_mmio_resp_bits_cmd,
  input  [63:0] io_mmio_resp_bits_rdata,
  output        io_frontend_req_ready,
  input         io_frontend_req_valid,
  input  [31:0] io_frontend_req_bits_addr,
  input  [2:0]  io_frontend_req_bits_size,
  input  [3:0]  io_frontend_req_bits_cmd,
  input  [7:0]  io_frontend_req_bits_wmask,
  input  [63:0] io_frontend_req_bits_wdata,
  input         io_frontend_resp_ready,
  output        io_frontend_resp_valid,
  output [3:0]  io_frontend_resp_bits_cmd,
  output [63:0] io_frontend_resp_bits_rdata,
  output [63:0] perfCnts_2,
  output [38:0] io_in_bits_decode_cf_pc,
  output [4:0]  io_wb_rfDest,
  input         io_extra_mtip,
  input         io_extra_meip_0,
  output        io_wb_rfWen,
  output [63:0] io_wb_rfData,
  input         io_extra_msip,
  output        io_in_valid_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [63:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [31:0] _RAND_22;
  reg [31:0] _RAND_23;
  reg [31:0] _RAND_24;
  reg [31:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [63:0] _RAND_28;
  reg [63:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [63:0] _RAND_31;
  reg [31:0] _RAND_32;
  reg [31:0] _RAND_33;
  reg [31:0] _RAND_34;
  reg [31:0] _RAND_35;
  reg [31:0] _RAND_36;
  reg [31:0] _RAND_37;
  reg [31:0] _RAND_38;
  reg [31:0] _RAND_39;
  reg [31:0] _RAND_40;
  reg [31:0] _RAND_41;
  reg [31:0] _RAND_42;
  reg [31:0] _RAND_43;
  reg [31:0] _RAND_44;
  reg [31:0] _RAND_45;
  reg [31:0] _RAND_46;
  reg [31:0] _RAND_47;
  reg [31:0] _RAND_48;
  reg [31:0] _RAND_49;
  reg [31:0] _RAND_50;
  reg [31:0] _RAND_51;
  reg [31:0] _RAND_52;
  reg [31:0] _RAND_53;
  reg [31:0] _RAND_54;
  reg [31:0] _RAND_55;
  reg [31:0] _RAND_56;
  reg [63:0] _RAND_57;
  reg [63:0] _RAND_58;
  reg [63:0] _RAND_59;
  reg [63:0] _RAND_60;
  reg [31:0] _RAND_61;
  reg [31:0] _RAND_62;
  reg [31:0] _RAND_63;
  reg [31:0] _RAND_64;
  reg [31:0] _RAND_65;
  reg [31:0] _RAND_66;
  reg [31:0] _RAND_67;
  reg [31:0] _RAND_68;
  reg [31:0] _RAND_69;
  reg [31:0] _RAND_70;
  reg [31:0] _RAND_71;
  reg [31:0] _RAND_72;
  reg [31:0] _RAND_73;
  reg [31:0] _RAND_74;
  reg [31:0] _RAND_75;
  reg [31:0] _RAND_76;
  reg [31:0] _RAND_77;
  reg [31:0] _RAND_78;
  reg [31:0] _RAND_79;
  reg [31:0] _RAND_80;
  reg [31:0] _RAND_81;
  reg [31:0] _RAND_82;
  reg [31:0] _RAND_83;
  reg [31:0] _RAND_84;
  reg [31:0] _RAND_85;
  reg [63:0] _RAND_86;
  reg [63:0] _RAND_87;
  reg [63:0] _RAND_88;
  reg [63:0] _RAND_89;
  reg [31:0] _RAND_90;
  reg [31:0] _RAND_91;
  reg [31:0] _RAND_92;
  reg [31:0] _RAND_93;
  reg [31:0] _RAND_94;
  reg [31:0] _RAND_95;
  reg [31:0] _RAND_96;
  reg [31:0] _RAND_97;
  reg [31:0] _RAND_98;
  reg [31:0] _RAND_99;
  reg [31:0] _RAND_100;
  reg [31:0] _RAND_101;
  reg [31:0] _RAND_102;
  reg [31:0] _RAND_103;
  reg [31:0] _RAND_104;
  reg [31:0] _RAND_105;
  reg [31:0] _RAND_106;
  reg [31:0] _RAND_107;
  reg [31:0] _RAND_108;
  reg [31:0] _RAND_109;
  reg [31:0] _RAND_110;
  reg [31:0] _RAND_111;
  reg [31:0] _RAND_112;
  reg [31:0] _RAND_113;
  reg [31:0] _RAND_114;
  reg [63:0] _RAND_115;
  reg [31:0] _RAND_116;
  reg [31:0] _RAND_117;
`endif // RANDOMIZE_REG_INIT
  wire  frontend_clock; // @[NutCore.scala 102:34]
  wire  frontend_reset; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_ready; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_valid; // @[NutCore.scala 102:34]
  wire [63:0] frontend_io_out_0_bits_cf_instr; // @[NutCore.scala 102:34]
  wire [38:0] frontend_io_out_0_bits_cf_pc; // @[NutCore.scala 102:34]
  wire [38:0] frontend_io_out_0_bits_cf_pnpc; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_exceptionVec_1; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_exceptionVec_2; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_exceptionVec_12; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_intrVec_0; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_intrVec_1; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_intrVec_2; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_intrVec_3; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_intrVec_4; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_intrVec_5; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_intrVec_6; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_intrVec_7; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_intrVec_8; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_intrVec_9; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_intrVec_10; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_intrVec_11; // @[NutCore.scala 102:34]
  wire [3:0] frontend_io_out_0_bits_cf_brIdx; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_cf_crossPageIPFFix; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_ctrl_src1Type; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_ctrl_src2Type; // @[NutCore.scala 102:34]
  wire [2:0] frontend_io_out_0_bits_ctrl_fuType; // @[NutCore.scala 102:34]
  wire [6:0] frontend_io_out_0_bits_ctrl_fuOpType; // @[NutCore.scala 102:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfSrc1; // @[NutCore.scala 102:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfSrc2; // @[NutCore.scala 102:34]
  wire  frontend_io_out_0_bits_ctrl_rfWen; // @[NutCore.scala 102:34]
  wire [4:0] frontend_io_out_0_bits_ctrl_rfDest; // @[NutCore.scala 102:34]
  wire [63:0] frontend_io_out_0_bits_data_imm; // @[NutCore.scala 102:34]
  wire  frontend_io_out_1_bits_cf_intrVec_0; // @[NutCore.scala 102:34]
  wire  frontend_io_out_1_bits_cf_intrVec_1; // @[NutCore.scala 102:34]
  wire  frontend_io_out_1_bits_cf_intrVec_2; // @[NutCore.scala 102:34]
  wire  frontend_io_out_1_bits_cf_intrVec_3; // @[NutCore.scala 102:34]
  wire  frontend_io_out_1_bits_cf_intrVec_4; // @[NutCore.scala 102:34]
  wire  frontend_io_out_1_bits_cf_intrVec_5; // @[NutCore.scala 102:34]
  wire  frontend_io_out_1_bits_cf_intrVec_6; // @[NutCore.scala 102:34]
  wire  frontend_io_out_1_bits_cf_intrVec_7; // @[NutCore.scala 102:34]
  wire  frontend_io_out_1_bits_cf_intrVec_8; // @[NutCore.scala 102:34]
  wire  frontend_io_out_1_bits_cf_intrVec_9; // @[NutCore.scala 102:34]
  wire  frontend_io_out_1_bits_cf_intrVec_10; // @[NutCore.scala 102:34]
  wire  frontend_io_out_1_bits_cf_intrVec_11; // @[NutCore.scala 102:34]
  wire  frontend_io_imem_req_ready; // @[NutCore.scala 102:34]
  wire  frontend_io_imem_req_valid; // @[NutCore.scala 102:34]
  wire [38:0] frontend_io_imem_req_bits_addr; // @[NutCore.scala 102:34]
  wire [86:0] frontend_io_imem_req_bits_user; // @[NutCore.scala 102:34]
  wire  frontend_io_imem_resp_ready; // @[NutCore.scala 102:34]
  wire  frontend_io_imem_resp_valid; // @[NutCore.scala 102:34]
  wire [63:0] frontend_io_imem_resp_bits_rdata; // @[NutCore.scala 102:34]
  wire [86:0] frontend_io_imem_resp_bits_user; // @[NutCore.scala 102:34]
  wire [3:0] frontend_io_flushVec; // @[NutCore.scala 102:34]
  wire  frontend_io_ipf; // @[NutCore.scala 102:34]
  wire [38:0] frontend_io_redirect_target; // @[NutCore.scala 102:34]
  wire  frontend_io_redirect_valid; // @[NutCore.scala 102:34]
  wire  frontend_flushICache; // @[NutCore.scala 102:34]
  wire  frontend__T_243_valid; // @[NutCore.scala 102:34]
  wire [38:0] frontend__T_243_pc; // @[NutCore.scala 102:34]
  wire  frontend__T_243_isMissPredict; // @[NutCore.scala 102:34]
  wire [38:0] frontend__T_243_actualTarget; // @[NutCore.scala 102:34]
  wire  frontend__T_243_actualTaken; // @[NutCore.scala 102:34]
  wire [6:0] frontend__T_243_fuOpType; // @[NutCore.scala 102:34]
  wire [1:0] frontend__T_243_btbType; // @[NutCore.scala 102:34]
  wire  frontend__T_243_isRVC; // @[NutCore.scala 102:34]
  wire  frontend_vmEnable; // @[NutCore.scala 102:34]
  wire [11:0] frontend_intrVec; // @[NutCore.scala 102:34]
  wire  frontend_flushTLB; // @[NutCore.scala 102:34]
  wire  Backend_inorder_clock; // @[NutCore.scala 144:25]
  wire  Backend_inorder_reset; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_ready; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_valid; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder_io_in_0_bits_cf_instr; // @[NutCore.scala 144:25]
  wire [38:0] Backend_inorder_io_in_0_bits_cf_pc; // @[NutCore.scala 144:25]
  wire [38:0] Backend_inorder_io_in_0_bits_cf_pnpc; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_exceptionVec_1; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_exceptionVec_2; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_exceptionVec_12; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_0; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_1; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_2; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_3; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_4; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_5; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_6; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_7; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_8; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_9; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_10; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_intrVec_11; // @[NutCore.scala 144:25]
  wire [3:0] Backend_inorder_io_in_0_bits_cf_brIdx; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_cf_crossPageIPFFix; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_ctrl_src1Type; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_ctrl_src2Type; // @[NutCore.scala 144:25]
  wire [2:0] Backend_inorder_io_in_0_bits_ctrl_fuType; // @[NutCore.scala 144:25]
  wire [6:0] Backend_inorder_io_in_0_bits_ctrl_fuOpType; // @[NutCore.scala 144:25]
  wire [4:0] Backend_inorder_io_in_0_bits_ctrl_rfSrc1; // @[NutCore.scala 144:25]
  wire [4:0] Backend_inorder_io_in_0_bits_ctrl_rfSrc2; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_0_bits_ctrl_rfWen; // @[NutCore.scala 144:25]
  wire [4:0] Backend_inorder_io_in_0_bits_ctrl_rfDest; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder_io_in_0_bits_data_imm; // @[NutCore.scala 144:25]
  wire [1:0] Backend_inorder_io_flush; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_dmem_req_ready; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_dmem_req_valid; // @[NutCore.scala 144:25]
  wire [38:0] Backend_inorder_io_dmem_req_bits_addr; // @[NutCore.scala 144:25]
  wire [2:0] Backend_inorder_io_dmem_req_bits_size; // @[NutCore.scala 144:25]
  wire [3:0] Backend_inorder_io_dmem_req_bits_cmd; // @[NutCore.scala 144:25]
  wire [7:0] Backend_inorder_io_dmem_req_bits_wmask; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder_io_dmem_req_bits_wdata; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_dmem_resp_valid; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder_io_dmem_resp_bits_rdata; // @[NutCore.scala 144:25]
  wire [1:0] Backend_inorder_io_memMMU_imem_priviledgeMode; // @[NutCore.scala 144:25]
  wire [1:0] Backend_inorder_io_memMMU_dmem_priviledgeMode; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_memMMU_dmem_status_sum; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_memMMU_dmem_status_mxr; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_memMMU_dmem_loadPF; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_memMMU_dmem_storePF; // @[NutCore.scala 144:25]
  wire [38:0] Backend_inorder_io_memMMU_dmem_addr; // @[NutCore.scala 144:25]
  wire [38:0] Backend_inorder_io_redirect_target; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_redirect_valid; // @[NutCore.scala 144:25]
  wire  Backend_inorder__T_38; // @[NutCore.scala 144:25]
  wire  Backend_inorder_flushICache; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder_perfCnts_2; // @[NutCore.scala 144:25]
  wire [38:0] Backend_inorder_io_in_bits_decode_cf_pc; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder_satp; // @[NutCore.scala 144:25]
  wire  Backend_inorder__T_243_valid; // @[NutCore.scala 144:25]
  wire [38:0] Backend_inorder__T_243_pc; // @[NutCore.scala 144:25]
  wire  Backend_inorder__T_243_isMissPredict; // @[NutCore.scala 144:25]
  wire [38:0] Backend_inorder__T_243_actualTarget; // @[NutCore.scala 144:25]
  wire  Backend_inorder__T_243_actualTaken; // @[NutCore.scala 144:25]
  wire [6:0] Backend_inorder__T_243_fuOpType; // @[NutCore.scala 144:25]
  wire [1:0] Backend_inorder__T_243_btbType; // @[NutCore.scala 144:25]
  wire  Backend_inorder__T_243_isRVC; // @[NutCore.scala 144:25]
  wire [4:0] Backend_inorder_io_wb_rfDest; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_extra_mtip; // @[NutCore.scala 144:25]
  wire  Backend_inorder_amoReq; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_extra_meip_0; // @[NutCore.scala 144:25]
  wire  Backend_inorder_vmEnable; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_wb_rfWen; // @[NutCore.scala 144:25]
  wire [63:0] Backend_inorder_io_wb_rfData; // @[NutCore.scala 144:25]
  wire [11:0] Backend_inorder_intrVec; // @[NutCore.scala 144:25]
  wire  Backend_inorder__T_37; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_extra_msip; // @[NutCore.scala 144:25]
  wire  Backend_inorder_flushTLB; // @[NutCore.scala 144:25]
  wire  Backend_inorder_io_in_valid_0; // @[NutCore.scala 144:25]
  wire  SimpleBusCrossbarNto1_clock; // @[NutCore.scala 148:26]
  wire  SimpleBusCrossbarNto1_reset; // @[NutCore.scala 148:26]
  wire  SimpleBusCrossbarNto1_io_in_0_req_ready; // @[NutCore.scala 148:26]
  wire  SimpleBusCrossbarNto1_io_in_0_req_valid; // @[NutCore.scala 148:26]
  wire [31:0] SimpleBusCrossbarNto1_io_in_0_req_bits_addr; // @[NutCore.scala 148:26]
  wire [3:0] SimpleBusCrossbarNto1_io_in_0_req_bits_cmd; // @[NutCore.scala 148:26]
  wire [7:0] SimpleBusCrossbarNto1_io_in_0_req_bits_wmask; // @[NutCore.scala 148:26]
  wire [63:0] SimpleBusCrossbarNto1_io_in_0_req_bits_wdata; // @[NutCore.scala 148:26]
  wire  SimpleBusCrossbarNto1_io_in_0_resp_valid; // @[NutCore.scala 148:26]
  wire [3:0] SimpleBusCrossbarNto1_io_in_0_resp_bits_cmd; // @[NutCore.scala 148:26]
  wire [63:0] SimpleBusCrossbarNto1_io_in_0_resp_bits_rdata; // @[NutCore.scala 148:26]
  wire  SimpleBusCrossbarNto1_io_in_1_req_ready; // @[NutCore.scala 148:26]
  wire  SimpleBusCrossbarNto1_io_in_1_req_valid; // @[NutCore.scala 148:26]
  wire [31:0] SimpleBusCrossbarNto1_io_in_1_req_bits_addr; // @[NutCore.scala 148:26]
  wire [2:0] SimpleBusCrossbarNto1_io_in_1_req_bits_size; // @[NutCore.scala 148:26]
  wire [3:0] SimpleBusCrossbarNto1_io_in_1_req_bits_cmd; // @[NutCore.scala 148:26]
  wire [7:0] SimpleBusCrossbarNto1_io_in_1_req_bits_wmask; // @[NutCore.scala 148:26]
  wire [63:0] SimpleBusCrossbarNto1_io_in_1_req_bits_wdata; // @[NutCore.scala 148:26]
  wire  SimpleBusCrossbarNto1_io_in_1_resp_valid; // @[NutCore.scala 148:26]
  wire [3:0] SimpleBusCrossbarNto1_io_in_1_resp_bits_cmd; // @[NutCore.scala 148:26]
  wire [63:0] SimpleBusCrossbarNto1_io_in_1_resp_bits_rdata; // @[NutCore.scala 148:26]
  wire  SimpleBusCrossbarNto1_io_out_req_ready; // @[NutCore.scala 148:26]
  wire  SimpleBusCrossbarNto1_io_out_req_valid; // @[NutCore.scala 148:26]
  wire [31:0] SimpleBusCrossbarNto1_io_out_req_bits_addr; // @[NutCore.scala 148:26]
  wire [2:0] SimpleBusCrossbarNto1_io_out_req_bits_size; // @[NutCore.scala 148:26]
  wire [3:0] SimpleBusCrossbarNto1_io_out_req_bits_cmd; // @[NutCore.scala 148:26]
  wire [7:0] SimpleBusCrossbarNto1_io_out_req_bits_wmask; // @[NutCore.scala 148:26]
  wire [63:0] SimpleBusCrossbarNto1_io_out_req_bits_wdata; // @[NutCore.scala 148:26]
  wire  SimpleBusCrossbarNto1_io_out_resp_ready; // @[NutCore.scala 148:26]
  wire  SimpleBusCrossbarNto1_io_out_resp_valid; // @[NutCore.scala 148:26]
  wire [3:0] SimpleBusCrossbarNto1_io_out_resp_bits_cmd; // @[NutCore.scala 148:26]
  wire [63:0] SimpleBusCrossbarNto1_io_out_resp_bits_rdata; // @[NutCore.scala 148:26]
  wire  SimpleBusCrossbarNto1_1_clock; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_reset; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_in_0_req_ready; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_in_0_req_valid; // @[NutCore.scala 149:26]
  wire [31:0] SimpleBusCrossbarNto1_1_io_in_0_req_bits_addr; // @[NutCore.scala 149:26]
  wire [2:0] SimpleBusCrossbarNto1_1_io_in_0_req_bits_size; // @[NutCore.scala 149:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_in_0_req_bits_cmd; // @[NutCore.scala 149:26]
  wire [7:0] SimpleBusCrossbarNto1_1_io_in_0_req_bits_wmask; // @[NutCore.scala 149:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_0_req_bits_wdata; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_in_0_resp_valid; // @[NutCore.scala 149:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_0_resp_bits_rdata; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_in_1_req_ready; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_in_1_req_valid; // @[NutCore.scala 149:26]
  wire [31:0] SimpleBusCrossbarNto1_1_io_in_1_req_bits_addr; // @[NutCore.scala 149:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_in_1_req_bits_cmd; // @[NutCore.scala 149:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_1_req_bits_wdata; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_in_1_resp_valid; // @[NutCore.scala 149:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_1_resp_bits_rdata; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_in_2_req_ready; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_in_2_req_valid; // @[NutCore.scala 149:26]
  wire [31:0] SimpleBusCrossbarNto1_1_io_in_2_req_bits_addr; // @[NutCore.scala 149:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_in_2_req_bits_cmd; // @[NutCore.scala 149:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_2_req_bits_wdata; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_in_2_resp_valid; // @[NutCore.scala 149:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_2_resp_bits_rdata; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_in_3_req_ready; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_in_3_req_valid; // @[NutCore.scala 149:26]
  wire [31:0] SimpleBusCrossbarNto1_1_io_in_3_req_bits_addr; // @[NutCore.scala 149:26]
  wire [2:0] SimpleBusCrossbarNto1_1_io_in_3_req_bits_size; // @[NutCore.scala 149:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_in_3_req_bits_cmd; // @[NutCore.scala 149:26]
  wire [7:0] SimpleBusCrossbarNto1_1_io_in_3_req_bits_wmask; // @[NutCore.scala 149:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_3_req_bits_wdata; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_in_3_resp_ready; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_in_3_resp_valid; // @[NutCore.scala 149:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_in_3_resp_bits_cmd; // @[NutCore.scala 149:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_in_3_resp_bits_rdata; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_out_req_ready; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_out_req_valid; // @[NutCore.scala 149:26]
  wire [31:0] SimpleBusCrossbarNto1_1_io_out_req_bits_addr; // @[NutCore.scala 149:26]
  wire [2:0] SimpleBusCrossbarNto1_1_io_out_req_bits_size; // @[NutCore.scala 149:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_out_req_bits_cmd; // @[NutCore.scala 149:26]
  wire [7:0] SimpleBusCrossbarNto1_1_io_out_req_bits_wmask; // @[NutCore.scala 149:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_out_req_bits_wdata; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_out_resp_ready; // @[NutCore.scala 149:26]
  wire  SimpleBusCrossbarNto1_1_io_out_resp_valid; // @[NutCore.scala 149:26]
  wire [3:0] SimpleBusCrossbarNto1_1_io_out_resp_bits_cmd; // @[NutCore.scala 149:26]
  wire [63:0] SimpleBusCrossbarNto1_1_io_out_resp_bits_rdata; // @[NutCore.scala 149:26]
  wire  EmbeddedTLB_clock; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_reset; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_in_req_ready; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_in_req_valid; // @[EmbeddedTLB.scala 427:23]
  wire [38:0] EmbeddedTLB_io_in_req_bits_addr; // @[EmbeddedTLB.scala 427:23]
  wire [86:0] EmbeddedTLB_io_in_req_bits_user; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_in_resp_ready; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_in_resp_valid; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_io_in_resp_bits_rdata; // @[EmbeddedTLB.scala 427:23]
  wire [86:0] EmbeddedTLB_io_in_resp_bits_user; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_out_req_ready; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_out_req_valid; // @[EmbeddedTLB.scala 427:23]
  wire [31:0] EmbeddedTLB_io_out_req_bits_addr; // @[EmbeddedTLB.scala 427:23]
  wire [86:0] EmbeddedTLB_io_out_req_bits_user; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_out_resp_ready; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_out_resp_valid; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_io_out_resp_bits_rdata; // @[EmbeddedTLB.scala 427:23]
  wire [86:0] EmbeddedTLB_io_out_resp_bits_user; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_mem_req_ready; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_mem_req_valid; // @[EmbeddedTLB.scala 427:23]
  wire [31:0] EmbeddedTLB_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 427:23]
  wire [3:0] EmbeddedTLB_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_mem_resp_valid; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_flush; // @[EmbeddedTLB.scala 427:23]
  wire [1:0] EmbeddedTLB_io_csrMMU_priviledgeMode; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_cacheEmpty; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_io_ipf; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_CSRSATP; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_MOUFlushTLB; // @[EmbeddedTLB.scala 427:23]
  wire  Cache_clock; // @[Cache.scala 678:35]
  wire  Cache_reset; // @[Cache.scala 678:35]
  wire  Cache_io_in_req_ready; // @[Cache.scala 678:35]
  wire  Cache_io_in_req_valid; // @[Cache.scala 678:35]
  wire [31:0] Cache_io_in_req_bits_addr; // @[Cache.scala 678:35]
  wire [86:0] Cache_io_in_req_bits_user; // @[Cache.scala 678:35]
  wire  Cache_io_in_resp_ready; // @[Cache.scala 678:35]
  wire  Cache_io_in_resp_valid; // @[Cache.scala 678:35]
  wire [63:0] Cache_io_in_resp_bits_rdata; // @[Cache.scala 678:35]
  wire [86:0] Cache_io_in_resp_bits_user; // @[Cache.scala 678:35]
  wire [1:0] Cache_io_flush; // @[Cache.scala 678:35]
  wire  Cache_io_out_mem_req_ready; // @[Cache.scala 678:35]
  wire  Cache_io_out_mem_req_valid; // @[Cache.scala 678:35]
  wire [31:0] Cache_io_out_mem_req_bits_addr; // @[Cache.scala 678:35]
  wire [3:0] Cache_io_out_mem_req_bits_cmd; // @[Cache.scala 678:35]
  wire [63:0] Cache_io_out_mem_req_bits_wdata; // @[Cache.scala 678:35]
  wire  Cache_io_out_mem_resp_valid; // @[Cache.scala 678:35]
  wire [3:0] Cache_io_out_mem_resp_bits_cmd; // @[Cache.scala 678:35]
  wire [63:0] Cache_io_out_mem_resp_bits_rdata; // @[Cache.scala 678:35]
  wire  Cache_io_mmio_req_ready; // @[Cache.scala 678:35]
  wire  Cache_io_mmio_req_valid; // @[Cache.scala 678:35]
  wire [31:0] Cache_io_mmio_req_bits_addr; // @[Cache.scala 678:35]
  wire  Cache_io_mmio_resp_valid; // @[Cache.scala 678:35]
  wire [63:0] Cache_io_mmio_resp_bits_rdata; // @[Cache.scala 678:35]
  wire  Cache_io_empty; // @[Cache.scala 678:35]
  wire  Cache_MOUFlushICache; // @[Cache.scala 678:35]
  wire  EmbeddedTLB_1_clock; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_reset; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_in_req_ready; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_in_req_valid; // @[EmbeddedTLB.scala 427:23]
  wire [38:0] EmbeddedTLB_1_io_in_req_bits_addr; // @[EmbeddedTLB.scala 427:23]
  wire [2:0] EmbeddedTLB_1_io_in_req_bits_size; // @[EmbeddedTLB.scala 427:23]
  wire [3:0] EmbeddedTLB_1_io_in_req_bits_cmd; // @[EmbeddedTLB.scala 427:23]
  wire [7:0] EmbeddedTLB_1_io_in_req_bits_wmask; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_1_io_in_req_bits_wdata; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_in_resp_valid; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_1_io_in_resp_bits_rdata; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_out_req_ready; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_out_req_valid; // @[EmbeddedTLB.scala 427:23]
  wire [31:0] EmbeddedTLB_1_io_out_req_bits_addr; // @[EmbeddedTLB.scala 427:23]
  wire [2:0] EmbeddedTLB_1_io_out_req_bits_size; // @[EmbeddedTLB.scala 427:23]
  wire [3:0] EmbeddedTLB_1_io_out_req_bits_cmd; // @[EmbeddedTLB.scala 427:23]
  wire [7:0] EmbeddedTLB_1_io_out_req_bits_wmask; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_1_io_out_req_bits_wdata; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_out_resp_valid; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_1_io_out_resp_bits_rdata; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_mem_req_ready; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_mem_req_valid; // @[EmbeddedTLB.scala 427:23]
  wire [31:0] EmbeddedTLB_1_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 427:23]
  wire [3:0] EmbeddedTLB_1_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_1_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_mem_resp_valid; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_1_io_mem_resp_bits_rdata; // @[EmbeddedTLB.scala 427:23]
  wire [1:0] EmbeddedTLB_1_io_csrMMU_priviledgeMode; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_csrMMU_status_sum; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_csrMMU_status_mxr; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_csrMMU_loadPF; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_io_csrMMU_storePF; // @[EmbeddedTLB.scala 427:23]
  wire [38:0] EmbeddedTLB_1_io_csrMMU_addr; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1__T_38_0; // @[EmbeddedTLB.scala 427:23]
  wire [63:0] EmbeddedTLB_1_CSRSATP; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_amoReq; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_vmEnable_0; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1__T_37_0; // @[EmbeddedTLB.scala 427:23]
  wire  EmbeddedTLB_1_MOUFlushTLB; // @[EmbeddedTLB.scala 427:23]
  wire  Cache_1_clock; // @[Cache.scala 678:35]
  wire  Cache_1_reset; // @[Cache.scala 678:35]
  wire  Cache_1_io_in_req_ready; // @[Cache.scala 678:35]
  wire  Cache_1_io_in_req_valid; // @[Cache.scala 678:35]
  wire [31:0] Cache_1_io_in_req_bits_addr; // @[Cache.scala 678:35]
  wire [2:0] Cache_1_io_in_req_bits_size; // @[Cache.scala 678:35]
  wire [3:0] Cache_1_io_in_req_bits_cmd; // @[Cache.scala 678:35]
  wire [7:0] Cache_1_io_in_req_bits_wmask; // @[Cache.scala 678:35]
  wire [63:0] Cache_1_io_in_req_bits_wdata; // @[Cache.scala 678:35]
  wire  Cache_1_io_in_resp_ready; // @[Cache.scala 678:35]
  wire  Cache_1_io_in_resp_valid; // @[Cache.scala 678:35]
  wire [3:0] Cache_1_io_in_resp_bits_cmd; // @[Cache.scala 678:35]
  wire [63:0] Cache_1_io_in_resp_bits_rdata; // @[Cache.scala 678:35]
  wire  Cache_1_io_out_mem_req_ready; // @[Cache.scala 678:35]
  wire  Cache_1_io_out_mem_req_valid; // @[Cache.scala 678:35]
  wire [31:0] Cache_1_io_out_mem_req_bits_addr; // @[Cache.scala 678:35]
  wire [3:0] Cache_1_io_out_mem_req_bits_cmd; // @[Cache.scala 678:35]
  wire [63:0] Cache_1_io_out_mem_req_bits_wdata; // @[Cache.scala 678:35]
  wire  Cache_1_io_out_mem_resp_valid; // @[Cache.scala 678:35]
  wire [3:0] Cache_1_io_out_mem_resp_bits_cmd; // @[Cache.scala 678:35]
  wire [63:0] Cache_1_io_out_mem_resp_bits_rdata; // @[Cache.scala 678:35]
  wire  Cache_1_io_out_coh_req_ready; // @[Cache.scala 678:35]
  wire  Cache_1_io_out_coh_req_valid; // @[Cache.scala 678:35]
  wire [31:0] Cache_1_io_out_coh_req_bits_addr; // @[Cache.scala 678:35]
  wire [63:0] Cache_1_io_out_coh_req_bits_wdata; // @[Cache.scala 678:35]
  wire  Cache_1_io_out_coh_resp_valid; // @[Cache.scala 678:35]
  wire [3:0] Cache_1_io_out_coh_resp_bits_cmd; // @[Cache.scala 678:35]
  wire [63:0] Cache_1_io_out_coh_resp_bits_rdata; // @[Cache.scala 678:35]
  wire  Cache_1_io_mmio_req_ready; // @[Cache.scala 678:35]
  wire  Cache_1_io_mmio_req_valid; // @[Cache.scala 678:35]
  wire [31:0] Cache_1_io_mmio_req_bits_addr; // @[Cache.scala 678:35]
  wire [2:0] Cache_1_io_mmio_req_bits_size; // @[Cache.scala 678:35]
  wire [3:0] Cache_1_io_mmio_req_bits_cmd; // @[Cache.scala 678:35]
  wire [7:0] Cache_1_io_mmio_req_bits_wmask; // @[Cache.scala 678:35]
  wire [63:0] Cache_1_io_mmio_req_bits_wdata; // @[Cache.scala 678:35]
  wire  Cache_1_io_mmio_resp_valid; // @[Cache.scala 678:35]
  wire [63:0] Cache_1_io_mmio_resp_bits_rdata; // @[Cache.scala 678:35]
  reg [63:0] _T_6_0_cf_instr; // @[PipelineVector.scala 29:29]
  reg [38:0] _T_6_0_cf_pc; // @[PipelineVector.scala 29:29]
  reg [38:0] _T_6_0_cf_pnpc; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_exceptionVec_1; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_exceptionVec_2; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_exceptionVec_12; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_intrVec_0; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_intrVec_1; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_intrVec_2; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_intrVec_3; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_intrVec_4; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_intrVec_5; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_intrVec_6; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_intrVec_7; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_intrVec_8; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_intrVec_9; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_intrVec_10; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_intrVec_11; // @[PipelineVector.scala 29:29]
  reg [3:0] _T_6_0_cf_brIdx; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_ctrl_src1Type; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_ctrl_src2Type; // @[PipelineVector.scala 29:29]
  reg [2:0] _T_6_0_ctrl_fuType; // @[PipelineVector.scala 29:29]
  reg [6:0] _T_6_0_ctrl_fuOpType; // @[PipelineVector.scala 29:29]
  reg [4:0] _T_6_0_ctrl_rfSrc1; // @[PipelineVector.scala 29:29]
  reg [4:0] _T_6_0_ctrl_rfSrc2; // @[PipelineVector.scala 29:29]
  reg  _T_6_0_ctrl_rfWen; // @[PipelineVector.scala 29:29]
  reg [4:0] _T_6_0_ctrl_rfDest; // @[PipelineVector.scala 29:29]
  reg [63:0] _T_6_0_data_imm; // @[PipelineVector.scala 29:29]
  reg [63:0] _T_6_1_cf_instr; // @[PipelineVector.scala 29:29]
  reg [38:0] _T_6_1_cf_pc; // @[PipelineVector.scala 29:29]
  reg [38:0] _T_6_1_cf_pnpc; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_exceptionVec_1; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_exceptionVec_2; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_exceptionVec_12; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_intrVec_0; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_intrVec_1; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_intrVec_2; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_intrVec_3; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_intrVec_4; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_intrVec_5; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_intrVec_6; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_intrVec_7; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_intrVec_8; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_intrVec_9; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_intrVec_10; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_intrVec_11; // @[PipelineVector.scala 29:29]
  reg [3:0] _T_6_1_cf_brIdx; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_ctrl_src1Type; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_ctrl_src2Type; // @[PipelineVector.scala 29:29]
  reg [2:0] _T_6_1_ctrl_fuType; // @[PipelineVector.scala 29:29]
  reg [6:0] _T_6_1_ctrl_fuOpType; // @[PipelineVector.scala 29:29]
  reg [4:0] _T_6_1_ctrl_rfSrc1; // @[PipelineVector.scala 29:29]
  reg [4:0] _T_6_1_ctrl_rfSrc2; // @[PipelineVector.scala 29:29]
  reg  _T_6_1_ctrl_rfWen; // @[PipelineVector.scala 29:29]
  reg [4:0] _T_6_1_ctrl_rfDest; // @[PipelineVector.scala 29:29]
  reg [63:0] _T_6_1_data_imm; // @[PipelineVector.scala 29:29]
  reg [63:0] _T_6_2_cf_instr; // @[PipelineVector.scala 29:29]
  reg [38:0] _T_6_2_cf_pc; // @[PipelineVector.scala 29:29]
  reg [38:0] _T_6_2_cf_pnpc; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_exceptionVec_1; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_exceptionVec_2; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_exceptionVec_12; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_intrVec_0; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_intrVec_1; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_intrVec_2; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_intrVec_3; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_intrVec_4; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_intrVec_5; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_intrVec_6; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_intrVec_7; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_intrVec_8; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_intrVec_9; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_intrVec_10; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_intrVec_11; // @[PipelineVector.scala 29:29]
  reg [3:0] _T_6_2_cf_brIdx; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_ctrl_src1Type; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_ctrl_src2Type; // @[PipelineVector.scala 29:29]
  reg [2:0] _T_6_2_ctrl_fuType; // @[PipelineVector.scala 29:29]
  reg [6:0] _T_6_2_ctrl_fuOpType; // @[PipelineVector.scala 29:29]
  reg [4:0] _T_6_2_ctrl_rfSrc1; // @[PipelineVector.scala 29:29]
  reg [4:0] _T_6_2_ctrl_rfSrc2; // @[PipelineVector.scala 29:29]
  reg  _T_6_2_ctrl_rfWen; // @[PipelineVector.scala 29:29]
  reg [4:0] _T_6_2_ctrl_rfDest; // @[PipelineVector.scala 29:29]
  reg [63:0] _T_6_2_data_imm; // @[PipelineVector.scala 29:29]
  reg [63:0] _T_6_3_cf_instr; // @[PipelineVector.scala 29:29]
  reg [38:0] _T_6_3_cf_pc; // @[PipelineVector.scala 29:29]
  reg [38:0] _T_6_3_cf_pnpc; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_exceptionVec_1; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_exceptionVec_2; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_exceptionVec_12; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_intrVec_0; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_intrVec_1; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_intrVec_2; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_intrVec_3; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_intrVec_4; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_intrVec_5; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_intrVec_6; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_intrVec_7; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_intrVec_8; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_intrVec_9; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_intrVec_10; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_intrVec_11; // @[PipelineVector.scala 29:29]
  reg [3:0] _T_6_3_cf_brIdx; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_cf_crossPageIPFFix; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_ctrl_src1Type; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_ctrl_src2Type; // @[PipelineVector.scala 29:29]
  reg [2:0] _T_6_3_ctrl_fuType; // @[PipelineVector.scala 29:29]
  reg [6:0] _T_6_3_ctrl_fuOpType; // @[PipelineVector.scala 29:29]
  reg [4:0] _T_6_3_ctrl_rfSrc1; // @[PipelineVector.scala 29:29]
  reg [4:0] _T_6_3_ctrl_rfSrc2; // @[PipelineVector.scala 29:29]
  reg  _T_6_3_ctrl_rfWen; // @[PipelineVector.scala 29:29]
  reg [4:0] _T_6_3_ctrl_rfDest; // @[PipelineVector.scala 29:29]
  reg [63:0] _T_6_3_data_imm; // @[PipelineVector.scala 29:29]
  reg [1:0] _T_7; // @[PipelineVector.scala 30:33]
  reg [1:0] _T_8; // @[PipelineVector.scala 31:33]
  wire [1:0] _T_11 = _T_7 + 2'h1; // @[PipelineVector.scala 33:63]
  wire  _T_12 = _T_11 != _T_8; // @[PipelineVector.scala 33:74]
  wire [1:0] _T_14 = _T_7 + 2'h2; // @[PipelineVector.scala 33:63]
  wire  _T_15 = _T_14 != _T_8; // @[PipelineVector.scala 33:74]
  wire  _T_17 = _T_12 & _T_15; // @[PipelineVector.scala 33:124]
  wire  _T_18_0 = frontend_io_out_0_valid; // @[PipelineVector.scala 36:27 PipelineVector.scala 37:20]
  wire [1:0] _T_19 = {{1'd0}, _T_18_0}; // @[PipelineVector.scala 40:46]
  wire  _T_20 = _T_19 >= 2'h1; // @[PipelineVector.scala 41:53]
  wire  _T_21 = _T_19 >= 2'h2; // @[PipelineVector.scala 41:53]
  wire  _T_22 = frontend_io_out_0_ready & frontend_io_out_0_valid; // @[Decoupled.scala 40:37]
  wire [2:0] _T_25 = {{1'd0}, _T_7}; // @[PipelineVector.scala 45:45]
  wire [63:0] _T_27_cf_instr = _T_18_0 ? frontend_io_out_0_bits_cf_instr : 64'h0; // @[PipelineVector.scala 45:69]
  wire [38:0] _T_27_cf_pc = _T_18_0 ? frontend_io_out_0_bits_cf_pc : 39'h0; // @[PipelineVector.scala 45:69]
  wire [38:0] _T_27_cf_pnpc = _T_18_0 ? frontend_io_out_0_bits_cf_pnpc : 39'h0; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_exceptionVec_1 = _T_18_0 & frontend_io_out_0_bits_cf_exceptionVec_1; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_exceptionVec_2 = _T_18_0 & frontend_io_out_0_bits_cf_exceptionVec_2; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_exceptionVec_12 = _T_18_0 & frontend_io_out_0_bits_cf_exceptionVec_12; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_intrVec_0 = _T_18_0 ? frontend_io_out_0_bits_cf_intrVec_0 : frontend_io_out_1_bits_cf_intrVec_0; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_intrVec_1 = _T_18_0 ? frontend_io_out_0_bits_cf_intrVec_1 : frontend_io_out_1_bits_cf_intrVec_1; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_intrVec_2 = _T_18_0 ? frontend_io_out_0_bits_cf_intrVec_2 : frontend_io_out_1_bits_cf_intrVec_2; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_intrVec_3 = _T_18_0 ? frontend_io_out_0_bits_cf_intrVec_3 : frontend_io_out_1_bits_cf_intrVec_3; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_intrVec_4 = _T_18_0 ? frontend_io_out_0_bits_cf_intrVec_4 : frontend_io_out_1_bits_cf_intrVec_4; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_intrVec_5 = _T_18_0 ? frontend_io_out_0_bits_cf_intrVec_5 : frontend_io_out_1_bits_cf_intrVec_5; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_intrVec_6 = _T_18_0 ? frontend_io_out_0_bits_cf_intrVec_6 : frontend_io_out_1_bits_cf_intrVec_6; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_intrVec_7 = _T_18_0 ? frontend_io_out_0_bits_cf_intrVec_7 : frontend_io_out_1_bits_cf_intrVec_7; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_intrVec_8 = _T_18_0 ? frontend_io_out_0_bits_cf_intrVec_8 : frontend_io_out_1_bits_cf_intrVec_8; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_intrVec_9 = _T_18_0 ? frontend_io_out_0_bits_cf_intrVec_9 : frontend_io_out_1_bits_cf_intrVec_9; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_intrVec_10 = _T_18_0 ? frontend_io_out_0_bits_cf_intrVec_10 : frontend_io_out_1_bits_cf_intrVec_10; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_intrVec_11 = _T_18_0 ? frontend_io_out_0_bits_cf_intrVec_11 : frontend_io_out_1_bits_cf_intrVec_11; // @[PipelineVector.scala 45:69]
  wire [3:0] _T_27_cf_brIdx = _T_18_0 ? frontend_io_out_0_bits_cf_brIdx : 4'h0; // @[PipelineVector.scala 45:69]
  wire  _T_27_cf_crossPageIPFFix = _T_18_0 & frontend_io_out_0_bits_cf_crossPageIPFFix; // @[PipelineVector.scala 45:69]
  wire  _T_27_ctrl_src1Type = _T_18_0 ? frontend_io_out_0_bits_ctrl_src1Type : 1'h1; // @[PipelineVector.scala 45:69]
  wire  _T_27_ctrl_src2Type = _T_18_0 ? frontend_io_out_0_bits_ctrl_src2Type : 1'h1; // @[PipelineVector.scala 45:69]
  wire [2:0] _T_27_ctrl_fuType = _T_18_0 ? frontend_io_out_0_bits_ctrl_fuType : 3'h3; // @[PipelineVector.scala 45:69]
  wire [6:0] _T_27_ctrl_fuOpType = _T_18_0 ? frontend_io_out_0_bits_ctrl_fuOpType : 7'h0; // @[PipelineVector.scala 45:69]
  wire [4:0] _T_27_ctrl_rfSrc1 = _T_18_0 ? frontend_io_out_0_bits_ctrl_rfSrc1 : 5'h0; // @[PipelineVector.scala 45:69]
  wire [4:0] _T_27_ctrl_rfSrc2 = _T_18_0 ? frontend_io_out_0_bits_ctrl_rfSrc2 : 5'h0; // @[PipelineVector.scala 45:69]
  wire  _T_27_ctrl_rfWen = _T_18_0 & frontend_io_out_0_bits_ctrl_rfWen; // @[PipelineVector.scala 45:69]
  wire [4:0] _T_27_ctrl_rfDest = _T_18_0 ? frontend_io_out_0_bits_ctrl_rfDest : 5'h0; // @[PipelineVector.scala 45:69]
  wire [63:0] _T_27_data_imm = _T_18_0 ? frontend_io_out_0_bits_data_imm : 64'h0; // @[PipelineVector.scala 45:69]
  wire  _GEN_56 = 2'h0 == _T_25[1:0] ? _T_27_ctrl_src2Type : _T_6_0_ctrl_src2Type; // @[PipelineVector.scala 45:63]
  wire  _GEN_57 = 2'h1 == _T_25[1:0] ? _T_27_ctrl_src2Type : _T_6_1_ctrl_src2Type; // @[PipelineVector.scala 45:63]
  wire  _GEN_58 = 2'h2 == _T_25[1:0] ? _T_27_ctrl_src2Type : _T_6_2_ctrl_src2Type; // @[PipelineVector.scala 45:63]
  wire  _GEN_59 = 2'h3 == _T_25[1:0] ? _T_27_ctrl_src2Type : _T_6_3_ctrl_src2Type; // @[PipelineVector.scala 45:63]
  wire  _GEN_60 = 2'h0 == _T_25[1:0] ? _T_27_ctrl_src1Type : _T_6_0_ctrl_src1Type; // @[PipelineVector.scala 45:63]
  wire  _GEN_61 = 2'h1 == _T_25[1:0] ? _T_27_ctrl_src1Type : _T_6_1_ctrl_src1Type; // @[PipelineVector.scala 45:63]
  wire  _GEN_62 = 2'h2 == _T_25[1:0] ? _T_27_ctrl_src1Type : _T_6_2_ctrl_src1Type; // @[PipelineVector.scala 45:63]
  wire  _GEN_63 = 2'h3 == _T_25[1:0] ? _T_27_ctrl_src1Type : _T_6_3_ctrl_src1Type; // @[PipelineVector.scala 45:63]
  wire  _GEN_268 = _T_20 ? _GEN_56 : _T_6_0_ctrl_src2Type; // @[PipelineVector.scala 45:29]
  wire  _GEN_269 = _T_20 ? _GEN_57 : _T_6_1_ctrl_src2Type; // @[PipelineVector.scala 45:29]
  wire  _GEN_270 = _T_20 ? _GEN_58 : _T_6_2_ctrl_src2Type; // @[PipelineVector.scala 45:29]
  wire  _GEN_271 = _T_20 ? _GEN_59 : _T_6_3_ctrl_src2Type; // @[PipelineVector.scala 45:29]
  wire  _GEN_272 = _T_20 ? _GEN_60 : _T_6_0_ctrl_src1Type; // @[PipelineVector.scala 45:29]
  wire  _GEN_273 = _T_20 ? _GEN_61 : _T_6_1_ctrl_src1Type; // @[PipelineVector.scala 45:29]
  wire  _GEN_274 = _T_20 ? _GEN_62 : _T_6_2_ctrl_src1Type; // @[PipelineVector.scala 45:29]
  wire  _GEN_275 = _T_20 ? _GEN_63 : _T_6_3_ctrl_src1Type; // @[PipelineVector.scala 45:29]
  wire [1:0] _T_29 = 2'h1 + _T_7; // @[PipelineVector.scala 46:45]
  wire  _GEN_1488 = 2'h0 == _T_29; // @[PipelineVector.scala 46:63]
  wire  _GEN_480 = _GEN_1488 | _GEN_268; // @[PipelineVector.scala 46:63]
  wire  _GEN_1489 = 2'h1 == _T_29; // @[PipelineVector.scala 46:63]
  wire  _GEN_481 = _GEN_1489 | _GEN_269; // @[PipelineVector.scala 46:63]
  wire  _GEN_1490 = 2'h2 == _T_29; // @[PipelineVector.scala 46:63]
  wire  _GEN_482 = _GEN_1490 | _GEN_270; // @[PipelineVector.scala 46:63]
  wire  _GEN_1491 = 2'h3 == _T_29; // @[PipelineVector.scala 46:63]
  wire  _GEN_483 = _GEN_1491 | _GEN_271; // @[PipelineVector.scala 46:63]
  wire  _GEN_484 = _GEN_1488 | _GEN_272; // @[PipelineVector.scala 46:63]
  wire  _GEN_485 = _GEN_1489 | _GEN_273; // @[PipelineVector.scala 46:63]
  wire  _GEN_486 = _GEN_1490 | _GEN_274; // @[PipelineVector.scala 46:63]
  wire  _GEN_487 = _GEN_1491 | _GEN_275; // @[PipelineVector.scala 46:63]
  wire  _T_6_T_29_cf_intrVec_0 = frontend_io_out_1_bits_cf_intrVec_0; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire  _T_6_T_29_cf_intrVec_1 = frontend_io_out_1_bits_cf_intrVec_1; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire  _T_6_T_29_cf_intrVec_2 = frontend_io_out_1_bits_cf_intrVec_2; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire  _T_6_T_29_cf_intrVec_3 = frontend_io_out_1_bits_cf_intrVec_3; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire  _T_6_T_29_cf_intrVec_4 = frontend_io_out_1_bits_cf_intrVec_4; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire  _T_6_T_29_cf_intrVec_5 = frontend_io_out_1_bits_cf_intrVec_5; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire  _T_6_T_29_cf_intrVec_6 = frontend_io_out_1_bits_cf_intrVec_6; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire  _T_6_T_29_cf_intrVec_7 = frontend_io_out_1_bits_cf_intrVec_7; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire  _T_6_T_29_cf_intrVec_8 = frontend_io_out_1_bits_cf_intrVec_8; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire  _T_6_T_29_cf_intrVec_9 = frontend_io_out_1_bits_cf_intrVec_9; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire  _T_6_T_29_cf_intrVec_10 = frontend_io_out_1_bits_cf_intrVec_10; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire  _T_6_T_29_cf_intrVec_11 = frontend_io_out_1_bits_cf_intrVec_11; // @[PipelineVector.scala 46:63 PipelineVector.scala 46:63]
  wire [1:0] _T_31 = _T_7 + _T_19; // @[PipelineVector.scala 47:42]
  wire  _T_32 = ~frontend_io_out_0_valid; // @[PipelineVector.scala 50:39]
  wire [63:0] _GEN_1114 = 2'h1 == _T_8 ? _T_6_1_cf_instr : _T_6_0_cf_instr; // @[PipelineVector.scala 55:15]
  wire [38:0] _GEN_1115 = 2'h1 == _T_8 ? _T_6_1_cf_pc : _T_6_0_cf_pc; // @[PipelineVector.scala 55:15]
  wire [38:0] _GEN_1116 = 2'h1 == _T_8 ? _T_6_1_cf_pnpc : _T_6_0_cf_pnpc; // @[PipelineVector.scala 55:15]
  wire  _GEN_1121 = 2'h1 == _T_8 ? _T_6_1_cf_exceptionVec_1 : _T_6_0_cf_exceptionVec_1; // @[PipelineVector.scala 55:15]
  wire  _GEN_1122 = 2'h1 == _T_8 ? _T_6_1_cf_exceptionVec_2 : _T_6_0_cf_exceptionVec_2; // @[PipelineVector.scala 55:15]
  wire  _GEN_1132 = 2'h1 == _T_8 ? _T_6_1_cf_exceptionVec_12 : _T_6_0_cf_exceptionVec_12; // @[PipelineVector.scala 55:15]
  wire  _GEN_1136 = 2'h1 == _T_8 ? _T_6_1_cf_intrVec_0 : _T_6_0_cf_intrVec_0; // @[PipelineVector.scala 55:15]
  wire  _GEN_1137 = 2'h1 == _T_8 ? _T_6_1_cf_intrVec_1 : _T_6_0_cf_intrVec_1; // @[PipelineVector.scala 55:15]
  wire  _GEN_1138 = 2'h1 == _T_8 ? _T_6_1_cf_intrVec_2 : _T_6_0_cf_intrVec_2; // @[PipelineVector.scala 55:15]
  wire  _GEN_1139 = 2'h1 == _T_8 ? _T_6_1_cf_intrVec_3 : _T_6_0_cf_intrVec_3; // @[PipelineVector.scala 55:15]
  wire  _GEN_1140 = 2'h1 == _T_8 ? _T_6_1_cf_intrVec_4 : _T_6_0_cf_intrVec_4; // @[PipelineVector.scala 55:15]
  wire  _GEN_1141 = 2'h1 == _T_8 ? _T_6_1_cf_intrVec_5 : _T_6_0_cf_intrVec_5; // @[PipelineVector.scala 55:15]
  wire  _GEN_1142 = 2'h1 == _T_8 ? _T_6_1_cf_intrVec_6 : _T_6_0_cf_intrVec_6; // @[PipelineVector.scala 55:15]
  wire  _GEN_1143 = 2'h1 == _T_8 ? _T_6_1_cf_intrVec_7 : _T_6_0_cf_intrVec_7; // @[PipelineVector.scala 55:15]
  wire  _GEN_1144 = 2'h1 == _T_8 ? _T_6_1_cf_intrVec_8 : _T_6_0_cf_intrVec_8; // @[PipelineVector.scala 55:15]
  wire  _GEN_1145 = 2'h1 == _T_8 ? _T_6_1_cf_intrVec_9 : _T_6_0_cf_intrVec_9; // @[PipelineVector.scala 55:15]
  wire  _GEN_1146 = 2'h1 == _T_8 ? _T_6_1_cf_intrVec_10 : _T_6_0_cf_intrVec_10; // @[PipelineVector.scala 55:15]
  wire  _GEN_1147 = 2'h1 == _T_8 ? _T_6_1_cf_intrVec_11 : _T_6_0_cf_intrVec_11; // @[PipelineVector.scala 55:15]
  wire [3:0] _GEN_1148 = 2'h1 == _T_8 ? _T_6_1_cf_brIdx : _T_6_0_cf_brIdx; // @[PipelineVector.scala 55:15]
  wire  _GEN_1150 = 2'h1 == _T_8 ? _T_6_1_cf_crossPageIPFFix : _T_6_0_cf_crossPageIPFFix; // @[PipelineVector.scala 55:15]
  wire  _GEN_1151 = 2'h1 == _T_8 ? _T_6_1_ctrl_src1Type : _T_6_0_ctrl_src1Type; // @[PipelineVector.scala 55:15]
  wire  _GEN_1152 = 2'h1 == _T_8 ? _T_6_1_ctrl_src2Type : _T_6_0_ctrl_src2Type; // @[PipelineVector.scala 55:15]
  wire [2:0] _GEN_1153 = 2'h1 == _T_8 ? _T_6_1_ctrl_fuType : _T_6_0_ctrl_fuType; // @[PipelineVector.scala 55:15]
  wire [6:0] _GEN_1154 = 2'h1 == _T_8 ? _T_6_1_ctrl_fuOpType : _T_6_0_ctrl_fuOpType; // @[PipelineVector.scala 55:15]
  wire [4:0] _GEN_1155 = 2'h1 == _T_8 ? _T_6_1_ctrl_rfSrc1 : _T_6_0_ctrl_rfSrc1; // @[PipelineVector.scala 55:15]
  wire [4:0] _GEN_1156 = 2'h1 == _T_8 ? _T_6_1_ctrl_rfSrc2 : _T_6_0_ctrl_rfSrc2; // @[PipelineVector.scala 55:15]
  wire  _GEN_1157 = 2'h1 == _T_8 ? _T_6_1_ctrl_rfWen : _T_6_0_ctrl_rfWen; // @[PipelineVector.scala 55:15]
  wire [4:0] _GEN_1158 = 2'h1 == _T_8 ? _T_6_1_ctrl_rfDest : _T_6_0_ctrl_rfDest; // @[PipelineVector.scala 55:15]
  wire [63:0] _GEN_1166 = 2'h1 == _T_8 ? _T_6_1_data_imm : _T_6_0_data_imm; // @[PipelineVector.scala 55:15]
  wire [63:0] _GEN_1167 = 2'h2 == _T_8 ? _T_6_2_cf_instr : _GEN_1114; // @[PipelineVector.scala 55:15]
  wire [38:0] _GEN_1168 = 2'h2 == _T_8 ? _T_6_2_cf_pc : _GEN_1115; // @[PipelineVector.scala 55:15]
  wire [38:0] _GEN_1169 = 2'h2 == _T_8 ? _T_6_2_cf_pnpc : _GEN_1116; // @[PipelineVector.scala 55:15]
  wire  _GEN_1174 = 2'h2 == _T_8 ? _T_6_2_cf_exceptionVec_1 : _GEN_1121; // @[PipelineVector.scala 55:15]
  wire  _GEN_1175 = 2'h2 == _T_8 ? _T_6_2_cf_exceptionVec_2 : _GEN_1122; // @[PipelineVector.scala 55:15]
  wire  _GEN_1185 = 2'h2 == _T_8 ? _T_6_2_cf_exceptionVec_12 : _GEN_1132; // @[PipelineVector.scala 55:15]
  wire  _GEN_1189 = 2'h2 == _T_8 ? _T_6_2_cf_intrVec_0 : _GEN_1136; // @[PipelineVector.scala 55:15]
  wire  _GEN_1190 = 2'h2 == _T_8 ? _T_6_2_cf_intrVec_1 : _GEN_1137; // @[PipelineVector.scala 55:15]
  wire  _GEN_1191 = 2'h2 == _T_8 ? _T_6_2_cf_intrVec_2 : _GEN_1138; // @[PipelineVector.scala 55:15]
  wire  _GEN_1192 = 2'h2 == _T_8 ? _T_6_2_cf_intrVec_3 : _GEN_1139; // @[PipelineVector.scala 55:15]
  wire  _GEN_1193 = 2'h2 == _T_8 ? _T_6_2_cf_intrVec_4 : _GEN_1140; // @[PipelineVector.scala 55:15]
  wire  _GEN_1194 = 2'h2 == _T_8 ? _T_6_2_cf_intrVec_5 : _GEN_1141; // @[PipelineVector.scala 55:15]
  wire  _GEN_1195 = 2'h2 == _T_8 ? _T_6_2_cf_intrVec_6 : _GEN_1142; // @[PipelineVector.scala 55:15]
  wire  _GEN_1196 = 2'h2 == _T_8 ? _T_6_2_cf_intrVec_7 : _GEN_1143; // @[PipelineVector.scala 55:15]
  wire  _GEN_1197 = 2'h2 == _T_8 ? _T_6_2_cf_intrVec_8 : _GEN_1144; // @[PipelineVector.scala 55:15]
  wire  _GEN_1198 = 2'h2 == _T_8 ? _T_6_2_cf_intrVec_9 : _GEN_1145; // @[PipelineVector.scala 55:15]
  wire  _GEN_1199 = 2'h2 == _T_8 ? _T_6_2_cf_intrVec_10 : _GEN_1146; // @[PipelineVector.scala 55:15]
  wire  _GEN_1200 = 2'h2 == _T_8 ? _T_6_2_cf_intrVec_11 : _GEN_1147; // @[PipelineVector.scala 55:15]
  wire [3:0] _GEN_1201 = 2'h2 == _T_8 ? _T_6_2_cf_brIdx : _GEN_1148; // @[PipelineVector.scala 55:15]
  wire  _GEN_1203 = 2'h2 == _T_8 ? _T_6_2_cf_crossPageIPFFix : _GEN_1150; // @[PipelineVector.scala 55:15]
  wire  _GEN_1204 = 2'h2 == _T_8 ? _T_6_2_ctrl_src1Type : _GEN_1151; // @[PipelineVector.scala 55:15]
  wire  _GEN_1205 = 2'h2 == _T_8 ? _T_6_2_ctrl_src2Type : _GEN_1152; // @[PipelineVector.scala 55:15]
  wire [2:0] _GEN_1206 = 2'h2 == _T_8 ? _T_6_2_ctrl_fuType : _GEN_1153; // @[PipelineVector.scala 55:15]
  wire [6:0] _GEN_1207 = 2'h2 == _T_8 ? _T_6_2_ctrl_fuOpType : _GEN_1154; // @[PipelineVector.scala 55:15]
  wire [4:0] _GEN_1208 = 2'h2 == _T_8 ? _T_6_2_ctrl_rfSrc1 : _GEN_1155; // @[PipelineVector.scala 55:15]
  wire [4:0] _GEN_1209 = 2'h2 == _T_8 ? _T_6_2_ctrl_rfSrc2 : _GEN_1156; // @[PipelineVector.scala 55:15]
  wire  _GEN_1210 = 2'h2 == _T_8 ? _T_6_2_ctrl_rfWen : _GEN_1157; // @[PipelineVector.scala 55:15]
  wire [4:0] _GEN_1211 = 2'h2 == _T_8 ? _T_6_2_ctrl_rfDest : _GEN_1158; // @[PipelineVector.scala 55:15]
  wire [63:0] _GEN_1219 = 2'h2 == _T_8 ? _T_6_2_data_imm : _GEN_1166; // @[PipelineVector.scala 55:15]
  wire  _T_41 = Backend_inorder_io_in_0_ready & Backend_inorder_io_in_0_valid; // @[Decoupled.scala 40:37]
  wire [1:0] _T_43 = {{1'd0}, _T_41}; // @[PipelineVector.scala 64:44]
  wire  _T_44 = _T_43 > 2'h0; // @[PipelineVector.scala 65:35]
  wire [1:0] _T_46 = _T_8 + _T_43; // @[PipelineVector.scala 67:42]
  Frontend_inorder frontend ( // @[NutCore.scala 102:34]
    .clock(frontend_clock),
    .reset(frontend_reset),
    .io_out_0_ready(frontend_io_out_0_ready),
    .io_out_0_valid(frontend_io_out_0_valid),
    .io_out_0_bits_cf_instr(frontend_io_out_0_bits_cf_instr),
    .io_out_0_bits_cf_pc(frontend_io_out_0_bits_cf_pc),
    .io_out_0_bits_cf_pnpc(frontend_io_out_0_bits_cf_pnpc),
    .io_out_0_bits_cf_exceptionVec_1(frontend_io_out_0_bits_cf_exceptionVec_1),
    .io_out_0_bits_cf_exceptionVec_2(frontend_io_out_0_bits_cf_exceptionVec_2),
    .io_out_0_bits_cf_exceptionVec_12(frontend_io_out_0_bits_cf_exceptionVec_12),
    .io_out_0_bits_cf_intrVec_0(frontend_io_out_0_bits_cf_intrVec_0),
    .io_out_0_bits_cf_intrVec_1(frontend_io_out_0_bits_cf_intrVec_1),
    .io_out_0_bits_cf_intrVec_2(frontend_io_out_0_bits_cf_intrVec_2),
    .io_out_0_bits_cf_intrVec_3(frontend_io_out_0_bits_cf_intrVec_3),
    .io_out_0_bits_cf_intrVec_4(frontend_io_out_0_bits_cf_intrVec_4),
    .io_out_0_bits_cf_intrVec_5(frontend_io_out_0_bits_cf_intrVec_5),
    .io_out_0_bits_cf_intrVec_6(frontend_io_out_0_bits_cf_intrVec_6),
    .io_out_0_bits_cf_intrVec_7(frontend_io_out_0_bits_cf_intrVec_7),
    .io_out_0_bits_cf_intrVec_8(frontend_io_out_0_bits_cf_intrVec_8),
    .io_out_0_bits_cf_intrVec_9(frontend_io_out_0_bits_cf_intrVec_9),
    .io_out_0_bits_cf_intrVec_10(frontend_io_out_0_bits_cf_intrVec_10),
    .io_out_0_bits_cf_intrVec_11(frontend_io_out_0_bits_cf_intrVec_11),
    .io_out_0_bits_cf_brIdx(frontend_io_out_0_bits_cf_brIdx),
    .io_out_0_bits_cf_crossPageIPFFix(frontend_io_out_0_bits_cf_crossPageIPFFix),
    .io_out_0_bits_ctrl_src1Type(frontend_io_out_0_bits_ctrl_src1Type),
    .io_out_0_bits_ctrl_src2Type(frontend_io_out_0_bits_ctrl_src2Type),
    .io_out_0_bits_ctrl_fuType(frontend_io_out_0_bits_ctrl_fuType),
    .io_out_0_bits_ctrl_fuOpType(frontend_io_out_0_bits_ctrl_fuOpType),
    .io_out_0_bits_ctrl_rfSrc1(frontend_io_out_0_bits_ctrl_rfSrc1),
    .io_out_0_bits_ctrl_rfSrc2(frontend_io_out_0_bits_ctrl_rfSrc2),
    .io_out_0_bits_ctrl_rfWen(frontend_io_out_0_bits_ctrl_rfWen),
    .io_out_0_bits_ctrl_rfDest(frontend_io_out_0_bits_ctrl_rfDest),
    .io_out_0_bits_data_imm(frontend_io_out_0_bits_data_imm),
    .io_out_1_bits_cf_intrVec_0(frontend_io_out_1_bits_cf_intrVec_0),
    .io_out_1_bits_cf_intrVec_1(frontend_io_out_1_bits_cf_intrVec_1),
    .io_out_1_bits_cf_intrVec_2(frontend_io_out_1_bits_cf_intrVec_2),
    .io_out_1_bits_cf_intrVec_3(frontend_io_out_1_bits_cf_intrVec_3),
    .io_out_1_bits_cf_intrVec_4(frontend_io_out_1_bits_cf_intrVec_4),
    .io_out_1_bits_cf_intrVec_5(frontend_io_out_1_bits_cf_intrVec_5),
    .io_out_1_bits_cf_intrVec_6(frontend_io_out_1_bits_cf_intrVec_6),
    .io_out_1_bits_cf_intrVec_7(frontend_io_out_1_bits_cf_intrVec_7),
    .io_out_1_bits_cf_intrVec_8(frontend_io_out_1_bits_cf_intrVec_8),
    .io_out_1_bits_cf_intrVec_9(frontend_io_out_1_bits_cf_intrVec_9),
    .io_out_1_bits_cf_intrVec_10(frontend_io_out_1_bits_cf_intrVec_10),
    .io_out_1_bits_cf_intrVec_11(frontend_io_out_1_bits_cf_intrVec_11),
    .io_imem_req_ready(frontend_io_imem_req_ready),
    .io_imem_req_valid(frontend_io_imem_req_valid),
    .io_imem_req_bits_addr(frontend_io_imem_req_bits_addr),
    .io_imem_req_bits_user(frontend_io_imem_req_bits_user),
    .io_imem_resp_ready(frontend_io_imem_resp_ready),
    .io_imem_resp_valid(frontend_io_imem_resp_valid),
    .io_imem_resp_bits_rdata(frontend_io_imem_resp_bits_rdata),
    .io_imem_resp_bits_user(frontend_io_imem_resp_bits_user),
    .io_flushVec(frontend_io_flushVec),
    .io_ipf(frontend_io_ipf),
    .io_redirect_target(frontend_io_redirect_target),
    .io_redirect_valid(frontend_io_redirect_valid),
    .flushICache(frontend_flushICache),
    ._T_243_valid(frontend__T_243_valid),
    ._T_243_pc(frontend__T_243_pc),
    ._T_243_isMissPredict(frontend__T_243_isMissPredict),
    ._T_243_actualTarget(frontend__T_243_actualTarget),
    ._T_243_actualTaken(frontend__T_243_actualTaken),
    ._T_243_fuOpType(frontend__T_243_fuOpType),
    ._T_243_btbType(frontend__T_243_btbType),
    ._T_243_isRVC(frontend__T_243_isRVC),
    .vmEnable(frontend_vmEnable),
    .intrVec(frontend_intrVec),
    .flushTLB(frontend_flushTLB)
  );
  Backend_inorder Backend_inorder ( // @[NutCore.scala 144:25]
    .clock(Backend_inorder_clock),
    .reset(Backend_inorder_reset),
    .io_in_0_ready(Backend_inorder_io_in_0_ready),
    .io_in_0_valid(Backend_inorder_io_in_0_valid),
    .io_in_0_bits_cf_instr(Backend_inorder_io_in_0_bits_cf_instr),
    .io_in_0_bits_cf_pc(Backend_inorder_io_in_0_bits_cf_pc),
    .io_in_0_bits_cf_pnpc(Backend_inorder_io_in_0_bits_cf_pnpc),
    .io_in_0_bits_cf_exceptionVec_1(Backend_inorder_io_in_0_bits_cf_exceptionVec_1),
    .io_in_0_bits_cf_exceptionVec_2(Backend_inorder_io_in_0_bits_cf_exceptionVec_2),
    .io_in_0_bits_cf_exceptionVec_12(Backend_inorder_io_in_0_bits_cf_exceptionVec_12),
    .io_in_0_bits_cf_intrVec_0(Backend_inorder_io_in_0_bits_cf_intrVec_0),
    .io_in_0_bits_cf_intrVec_1(Backend_inorder_io_in_0_bits_cf_intrVec_1),
    .io_in_0_bits_cf_intrVec_2(Backend_inorder_io_in_0_bits_cf_intrVec_2),
    .io_in_0_bits_cf_intrVec_3(Backend_inorder_io_in_0_bits_cf_intrVec_3),
    .io_in_0_bits_cf_intrVec_4(Backend_inorder_io_in_0_bits_cf_intrVec_4),
    .io_in_0_bits_cf_intrVec_5(Backend_inorder_io_in_0_bits_cf_intrVec_5),
    .io_in_0_bits_cf_intrVec_6(Backend_inorder_io_in_0_bits_cf_intrVec_6),
    .io_in_0_bits_cf_intrVec_7(Backend_inorder_io_in_0_bits_cf_intrVec_7),
    .io_in_0_bits_cf_intrVec_8(Backend_inorder_io_in_0_bits_cf_intrVec_8),
    .io_in_0_bits_cf_intrVec_9(Backend_inorder_io_in_0_bits_cf_intrVec_9),
    .io_in_0_bits_cf_intrVec_10(Backend_inorder_io_in_0_bits_cf_intrVec_10),
    .io_in_0_bits_cf_intrVec_11(Backend_inorder_io_in_0_bits_cf_intrVec_11),
    .io_in_0_bits_cf_brIdx(Backend_inorder_io_in_0_bits_cf_brIdx),
    .io_in_0_bits_cf_crossPageIPFFix(Backend_inorder_io_in_0_bits_cf_crossPageIPFFix),
    .io_in_0_bits_ctrl_src1Type(Backend_inorder_io_in_0_bits_ctrl_src1Type),
    .io_in_0_bits_ctrl_src2Type(Backend_inorder_io_in_0_bits_ctrl_src2Type),
    .io_in_0_bits_ctrl_fuType(Backend_inorder_io_in_0_bits_ctrl_fuType),
    .io_in_0_bits_ctrl_fuOpType(Backend_inorder_io_in_0_bits_ctrl_fuOpType),
    .io_in_0_bits_ctrl_rfSrc1(Backend_inorder_io_in_0_bits_ctrl_rfSrc1),
    .io_in_0_bits_ctrl_rfSrc2(Backend_inorder_io_in_0_bits_ctrl_rfSrc2),
    .io_in_0_bits_ctrl_rfWen(Backend_inorder_io_in_0_bits_ctrl_rfWen),
    .io_in_0_bits_ctrl_rfDest(Backend_inorder_io_in_0_bits_ctrl_rfDest),
    .io_in_0_bits_data_imm(Backend_inorder_io_in_0_bits_data_imm),
    .io_flush(Backend_inorder_io_flush),
    .io_dmem_req_ready(Backend_inorder_io_dmem_req_ready),
    .io_dmem_req_valid(Backend_inorder_io_dmem_req_valid),
    .io_dmem_req_bits_addr(Backend_inorder_io_dmem_req_bits_addr),
    .io_dmem_req_bits_size(Backend_inorder_io_dmem_req_bits_size),
    .io_dmem_req_bits_cmd(Backend_inorder_io_dmem_req_bits_cmd),
    .io_dmem_req_bits_wmask(Backend_inorder_io_dmem_req_bits_wmask),
    .io_dmem_req_bits_wdata(Backend_inorder_io_dmem_req_bits_wdata),
    .io_dmem_resp_valid(Backend_inorder_io_dmem_resp_valid),
    .io_dmem_resp_bits_rdata(Backend_inorder_io_dmem_resp_bits_rdata),
    .io_memMMU_imem_priviledgeMode(Backend_inorder_io_memMMU_imem_priviledgeMode),
    .io_memMMU_dmem_priviledgeMode(Backend_inorder_io_memMMU_dmem_priviledgeMode),
    .io_memMMU_dmem_status_sum(Backend_inorder_io_memMMU_dmem_status_sum),
    .io_memMMU_dmem_status_mxr(Backend_inorder_io_memMMU_dmem_status_mxr),
    .io_memMMU_dmem_loadPF(Backend_inorder_io_memMMU_dmem_loadPF),
    .io_memMMU_dmem_storePF(Backend_inorder_io_memMMU_dmem_storePF),
    .io_memMMU_dmem_addr(Backend_inorder_io_memMMU_dmem_addr),
    .io_redirect_target(Backend_inorder_io_redirect_target),
    .io_redirect_valid(Backend_inorder_io_redirect_valid),
    ._T_38(Backend_inorder__T_38),
    .flushICache(Backend_inorder_flushICache),
    .perfCnts_2(Backend_inorder_perfCnts_2),
    .io_in_bits_decode_cf_pc(Backend_inorder_io_in_bits_decode_cf_pc),
    .satp(Backend_inorder_satp),
    ._T_243_valid(Backend_inorder__T_243_valid),
    ._T_243_pc(Backend_inorder__T_243_pc),
    ._T_243_isMissPredict(Backend_inorder__T_243_isMissPredict),
    ._T_243_actualTarget(Backend_inorder__T_243_actualTarget),
    ._T_243_actualTaken(Backend_inorder__T_243_actualTaken),
    ._T_243_fuOpType(Backend_inorder__T_243_fuOpType),
    ._T_243_btbType(Backend_inorder__T_243_btbType),
    ._T_243_isRVC(Backend_inorder__T_243_isRVC),
    .io_wb_rfDest(Backend_inorder_io_wb_rfDest),
    .io_extra_mtip(Backend_inorder_io_extra_mtip),
    .amoReq(Backend_inorder_amoReq),
    .io_extra_meip_0(Backend_inorder_io_extra_meip_0),
    .vmEnable(Backend_inorder_vmEnable),
    .io_wb_rfWen(Backend_inorder_io_wb_rfWen),
    .io_wb_rfData(Backend_inorder_io_wb_rfData),
    .intrVec(Backend_inorder_intrVec),
    ._T_37(Backend_inorder__T_37),
    .io_extra_msip(Backend_inorder_io_extra_msip),
    .flushTLB(Backend_inorder_flushTLB),
    .io_in_valid_0(Backend_inorder_io_in_valid_0)
  );
  SimpleBusCrossbarNto1 SimpleBusCrossbarNto1 ( // @[NutCore.scala 148:26]
    .clock(SimpleBusCrossbarNto1_clock),
    .reset(SimpleBusCrossbarNto1_reset),
    .io_in_0_req_ready(SimpleBusCrossbarNto1_io_in_0_req_ready),
    .io_in_0_req_valid(SimpleBusCrossbarNto1_io_in_0_req_valid),
    .io_in_0_req_bits_addr(SimpleBusCrossbarNto1_io_in_0_req_bits_addr),
    .io_in_0_req_bits_cmd(SimpleBusCrossbarNto1_io_in_0_req_bits_cmd),
    .io_in_0_req_bits_wmask(SimpleBusCrossbarNto1_io_in_0_req_bits_wmask),
    .io_in_0_req_bits_wdata(SimpleBusCrossbarNto1_io_in_0_req_bits_wdata),
    .io_in_0_resp_valid(SimpleBusCrossbarNto1_io_in_0_resp_valid),
    .io_in_0_resp_bits_cmd(SimpleBusCrossbarNto1_io_in_0_resp_bits_cmd),
    .io_in_0_resp_bits_rdata(SimpleBusCrossbarNto1_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(SimpleBusCrossbarNto1_io_in_1_req_ready),
    .io_in_1_req_valid(SimpleBusCrossbarNto1_io_in_1_req_valid),
    .io_in_1_req_bits_addr(SimpleBusCrossbarNto1_io_in_1_req_bits_addr),
    .io_in_1_req_bits_size(SimpleBusCrossbarNto1_io_in_1_req_bits_size),
    .io_in_1_req_bits_cmd(SimpleBusCrossbarNto1_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wmask(SimpleBusCrossbarNto1_io_in_1_req_bits_wmask),
    .io_in_1_req_bits_wdata(SimpleBusCrossbarNto1_io_in_1_req_bits_wdata),
    .io_in_1_resp_valid(SimpleBusCrossbarNto1_io_in_1_resp_valid),
    .io_in_1_resp_bits_cmd(SimpleBusCrossbarNto1_io_in_1_resp_bits_cmd),
    .io_in_1_resp_bits_rdata(SimpleBusCrossbarNto1_io_in_1_resp_bits_rdata),
    .io_out_req_ready(SimpleBusCrossbarNto1_io_out_req_ready),
    .io_out_req_valid(SimpleBusCrossbarNto1_io_out_req_valid),
    .io_out_req_bits_addr(SimpleBusCrossbarNto1_io_out_req_bits_addr),
    .io_out_req_bits_size(SimpleBusCrossbarNto1_io_out_req_bits_size),
    .io_out_req_bits_cmd(SimpleBusCrossbarNto1_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(SimpleBusCrossbarNto1_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(SimpleBusCrossbarNto1_io_out_req_bits_wdata),
    .io_out_resp_ready(SimpleBusCrossbarNto1_io_out_resp_ready),
    .io_out_resp_valid(SimpleBusCrossbarNto1_io_out_resp_valid),
    .io_out_resp_bits_cmd(SimpleBusCrossbarNto1_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(SimpleBusCrossbarNto1_io_out_resp_bits_rdata)
  );
  SimpleBusCrossbarNto1_1 SimpleBusCrossbarNto1_1 ( // @[NutCore.scala 149:26]
    .clock(SimpleBusCrossbarNto1_1_clock),
    .reset(SimpleBusCrossbarNto1_1_reset),
    .io_in_0_req_ready(SimpleBusCrossbarNto1_1_io_in_0_req_ready),
    .io_in_0_req_valid(SimpleBusCrossbarNto1_1_io_in_0_req_valid),
    .io_in_0_req_bits_addr(SimpleBusCrossbarNto1_1_io_in_0_req_bits_addr),
    .io_in_0_req_bits_size(SimpleBusCrossbarNto1_1_io_in_0_req_bits_size),
    .io_in_0_req_bits_cmd(SimpleBusCrossbarNto1_1_io_in_0_req_bits_cmd),
    .io_in_0_req_bits_wmask(SimpleBusCrossbarNto1_1_io_in_0_req_bits_wmask),
    .io_in_0_req_bits_wdata(SimpleBusCrossbarNto1_1_io_in_0_req_bits_wdata),
    .io_in_0_resp_valid(SimpleBusCrossbarNto1_1_io_in_0_resp_valid),
    .io_in_0_resp_bits_rdata(SimpleBusCrossbarNto1_1_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(SimpleBusCrossbarNto1_1_io_in_1_req_ready),
    .io_in_1_req_valid(SimpleBusCrossbarNto1_1_io_in_1_req_valid),
    .io_in_1_req_bits_addr(SimpleBusCrossbarNto1_1_io_in_1_req_bits_addr),
    .io_in_1_req_bits_cmd(SimpleBusCrossbarNto1_1_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wdata(SimpleBusCrossbarNto1_1_io_in_1_req_bits_wdata),
    .io_in_1_resp_valid(SimpleBusCrossbarNto1_1_io_in_1_resp_valid),
    .io_in_1_resp_bits_rdata(SimpleBusCrossbarNto1_1_io_in_1_resp_bits_rdata),
    .io_in_2_req_ready(SimpleBusCrossbarNto1_1_io_in_2_req_ready),
    .io_in_2_req_valid(SimpleBusCrossbarNto1_1_io_in_2_req_valid),
    .io_in_2_req_bits_addr(SimpleBusCrossbarNto1_1_io_in_2_req_bits_addr),
    .io_in_2_req_bits_cmd(SimpleBusCrossbarNto1_1_io_in_2_req_bits_cmd),
    .io_in_2_req_bits_wdata(SimpleBusCrossbarNto1_1_io_in_2_req_bits_wdata),
    .io_in_2_resp_valid(SimpleBusCrossbarNto1_1_io_in_2_resp_valid),
    .io_in_2_resp_bits_rdata(SimpleBusCrossbarNto1_1_io_in_2_resp_bits_rdata),
    .io_in_3_req_ready(SimpleBusCrossbarNto1_1_io_in_3_req_ready),
    .io_in_3_req_valid(SimpleBusCrossbarNto1_1_io_in_3_req_valid),
    .io_in_3_req_bits_addr(SimpleBusCrossbarNto1_1_io_in_3_req_bits_addr),
    .io_in_3_req_bits_size(SimpleBusCrossbarNto1_1_io_in_3_req_bits_size),
    .io_in_3_req_bits_cmd(SimpleBusCrossbarNto1_1_io_in_3_req_bits_cmd),
    .io_in_3_req_bits_wmask(SimpleBusCrossbarNto1_1_io_in_3_req_bits_wmask),
    .io_in_3_req_bits_wdata(SimpleBusCrossbarNto1_1_io_in_3_req_bits_wdata),
    .io_in_3_resp_ready(SimpleBusCrossbarNto1_1_io_in_3_resp_ready),
    .io_in_3_resp_valid(SimpleBusCrossbarNto1_1_io_in_3_resp_valid),
    .io_in_3_resp_bits_cmd(SimpleBusCrossbarNto1_1_io_in_3_resp_bits_cmd),
    .io_in_3_resp_bits_rdata(SimpleBusCrossbarNto1_1_io_in_3_resp_bits_rdata),
    .io_out_req_ready(SimpleBusCrossbarNto1_1_io_out_req_ready),
    .io_out_req_valid(SimpleBusCrossbarNto1_1_io_out_req_valid),
    .io_out_req_bits_addr(SimpleBusCrossbarNto1_1_io_out_req_bits_addr),
    .io_out_req_bits_size(SimpleBusCrossbarNto1_1_io_out_req_bits_size),
    .io_out_req_bits_cmd(SimpleBusCrossbarNto1_1_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(SimpleBusCrossbarNto1_1_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(SimpleBusCrossbarNto1_1_io_out_req_bits_wdata),
    .io_out_resp_ready(SimpleBusCrossbarNto1_1_io_out_resp_ready),
    .io_out_resp_valid(SimpleBusCrossbarNto1_1_io_out_resp_valid),
    .io_out_resp_bits_cmd(SimpleBusCrossbarNto1_1_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(SimpleBusCrossbarNto1_1_io_out_resp_bits_rdata)
  );
  EmbeddedTLB EmbeddedTLB ( // @[EmbeddedTLB.scala 427:23]
    .clock(EmbeddedTLB_clock),
    .reset(EmbeddedTLB_reset),
    .io_in_req_ready(EmbeddedTLB_io_in_req_ready),
    .io_in_req_valid(EmbeddedTLB_io_in_req_valid),
    .io_in_req_bits_addr(EmbeddedTLB_io_in_req_bits_addr),
    .io_in_req_bits_user(EmbeddedTLB_io_in_req_bits_user),
    .io_in_resp_ready(EmbeddedTLB_io_in_resp_ready),
    .io_in_resp_valid(EmbeddedTLB_io_in_resp_valid),
    .io_in_resp_bits_rdata(EmbeddedTLB_io_in_resp_bits_rdata),
    .io_in_resp_bits_user(EmbeddedTLB_io_in_resp_bits_user),
    .io_out_req_ready(EmbeddedTLB_io_out_req_ready),
    .io_out_req_valid(EmbeddedTLB_io_out_req_valid),
    .io_out_req_bits_addr(EmbeddedTLB_io_out_req_bits_addr),
    .io_out_req_bits_user(EmbeddedTLB_io_out_req_bits_user),
    .io_out_resp_ready(EmbeddedTLB_io_out_resp_ready),
    .io_out_resp_valid(EmbeddedTLB_io_out_resp_valid),
    .io_out_resp_bits_rdata(EmbeddedTLB_io_out_resp_bits_rdata),
    .io_out_resp_bits_user(EmbeddedTLB_io_out_resp_bits_user),
    .io_mem_req_ready(EmbeddedTLB_io_mem_req_ready),
    .io_mem_req_valid(EmbeddedTLB_io_mem_req_valid),
    .io_mem_req_bits_addr(EmbeddedTLB_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(EmbeddedTLB_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(EmbeddedTLB_io_mem_req_bits_wdata),
    .io_mem_resp_valid(EmbeddedTLB_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(EmbeddedTLB_io_mem_resp_bits_rdata),
    .io_flush(EmbeddedTLB_io_flush),
    .io_csrMMU_priviledgeMode(EmbeddedTLB_io_csrMMU_priviledgeMode),
    .io_cacheEmpty(EmbeddedTLB_io_cacheEmpty),
    .io_ipf(EmbeddedTLB_io_ipf),
    .CSRSATP(EmbeddedTLB_CSRSATP),
    .MOUFlushTLB(EmbeddedTLB_MOUFlushTLB)
  );
  Cache Cache ( // @[Cache.scala 678:35]
    .clock(Cache_clock),
    .reset(Cache_reset),
    .io_in_req_ready(Cache_io_in_req_ready),
    .io_in_req_valid(Cache_io_in_req_valid),
    .io_in_req_bits_addr(Cache_io_in_req_bits_addr),
    .io_in_req_bits_user(Cache_io_in_req_bits_user),
    .io_in_resp_ready(Cache_io_in_resp_ready),
    .io_in_resp_valid(Cache_io_in_resp_valid),
    .io_in_resp_bits_rdata(Cache_io_in_resp_bits_rdata),
    .io_in_resp_bits_user(Cache_io_in_resp_bits_user),
    .io_flush(Cache_io_flush),
    .io_out_mem_req_ready(Cache_io_out_mem_req_ready),
    .io_out_mem_req_valid(Cache_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(Cache_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_cmd(Cache_io_out_mem_req_bits_cmd),
    .io_out_mem_req_bits_wdata(Cache_io_out_mem_req_bits_wdata),
    .io_out_mem_resp_valid(Cache_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(Cache_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(Cache_io_out_mem_resp_bits_rdata),
    .io_mmio_req_ready(Cache_io_mmio_req_ready),
    .io_mmio_req_valid(Cache_io_mmio_req_valid),
    .io_mmio_req_bits_addr(Cache_io_mmio_req_bits_addr),
    .io_mmio_resp_valid(Cache_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(Cache_io_mmio_resp_bits_rdata),
    .io_empty(Cache_io_empty),
    .MOUFlushICache(Cache_MOUFlushICache)
  );
  EmbeddedTLB_1 EmbeddedTLB_1 ( // @[EmbeddedTLB.scala 427:23]
    .clock(EmbeddedTLB_1_clock),
    .reset(EmbeddedTLB_1_reset),
    .io_in_req_ready(EmbeddedTLB_1_io_in_req_ready),
    .io_in_req_valid(EmbeddedTLB_1_io_in_req_valid),
    .io_in_req_bits_addr(EmbeddedTLB_1_io_in_req_bits_addr),
    .io_in_req_bits_size(EmbeddedTLB_1_io_in_req_bits_size),
    .io_in_req_bits_cmd(EmbeddedTLB_1_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(EmbeddedTLB_1_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(EmbeddedTLB_1_io_in_req_bits_wdata),
    .io_in_resp_valid(EmbeddedTLB_1_io_in_resp_valid),
    .io_in_resp_bits_rdata(EmbeddedTLB_1_io_in_resp_bits_rdata),
    .io_out_req_ready(EmbeddedTLB_1_io_out_req_ready),
    .io_out_req_valid(EmbeddedTLB_1_io_out_req_valid),
    .io_out_req_bits_addr(EmbeddedTLB_1_io_out_req_bits_addr),
    .io_out_req_bits_size(EmbeddedTLB_1_io_out_req_bits_size),
    .io_out_req_bits_cmd(EmbeddedTLB_1_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(EmbeddedTLB_1_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(EmbeddedTLB_1_io_out_req_bits_wdata),
    .io_out_resp_valid(EmbeddedTLB_1_io_out_resp_valid),
    .io_out_resp_bits_rdata(EmbeddedTLB_1_io_out_resp_bits_rdata),
    .io_mem_req_ready(EmbeddedTLB_1_io_mem_req_ready),
    .io_mem_req_valid(EmbeddedTLB_1_io_mem_req_valid),
    .io_mem_req_bits_addr(EmbeddedTLB_1_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(EmbeddedTLB_1_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(EmbeddedTLB_1_io_mem_req_bits_wdata),
    .io_mem_resp_valid(EmbeddedTLB_1_io_mem_resp_valid),
    .io_mem_resp_bits_rdata(EmbeddedTLB_1_io_mem_resp_bits_rdata),
    .io_csrMMU_priviledgeMode(EmbeddedTLB_1_io_csrMMU_priviledgeMode),
    .io_csrMMU_status_sum(EmbeddedTLB_1_io_csrMMU_status_sum),
    .io_csrMMU_status_mxr(EmbeddedTLB_1_io_csrMMU_status_mxr),
    .io_csrMMU_loadPF(EmbeddedTLB_1_io_csrMMU_loadPF),
    .io_csrMMU_storePF(EmbeddedTLB_1_io_csrMMU_storePF),
    .io_csrMMU_addr(EmbeddedTLB_1_io_csrMMU_addr),
    ._T_38_0(EmbeddedTLB_1__T_38_0),
    .CSRSATP(EmbeddedTLB_1_CSRSATP),
    .amoReq(EmbeddedTLB_1_amoReq),
    .vmEnable_0(EmbeddedTLB_1_vmEnable_0),
    ._T_37_0(EmbeddedTLB_1__T_37_0),
    .MOUFlushTLB(EmbeddedTLB_1_MOUFlushTLB)
  );
  Cache_1 Cache_1 ( // @[Cache.scala 678:35]
    .clock(Cache_1_clock),
    .reset(Cache_1_reset),
    .io_in_req_ready(Cache_1_io_in_req_ready),
    .io_in_req_valid(Cache_1_io_in_req_valid),
    .io_in_req_bits_addr(Cache_1_io_in_req_bits_addr),
    .io_in_req_bits_size(Cache_1_io_in_req_bits_size),
    .io_in_req_bits_cmd(Cache_1_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(Cache_1_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(Cache_1_io_in_req_bits_wdata),
    .io_in_resp_ready(Cache_1_io_in_resp_ready),
    .io_in_resp_valid(Cache_1_io_in_resp_valid),
    .io_in_resp_bits_cmd(Cache_1_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(Cache_1_io_in_resp_bits_rdata),
    .io_out_mem_req_ready(Cache_1_io_out_mem_req_ready),
    .io_out_mem_req_valid(Cache_1_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(Cache_1_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_cmd(Cache_1_io_out_mem_req_bits_cmd),
    .io_out_mem_req_bits_wdata(Cache_1_io_out_mem_req_bits_wdata),
    .io_out_mem_resp_valid(Cache_1_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(Cache_1_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(Cache_1_io_out_mem_resp_bits_rdata),
    .io_out_coh_req_ready(Cache_1_io_out_coh_req_ready),
    .io_out_coh_req_valid(Cache_1_io_out_coh_req_valid),
    .io_out_coh_req_bits_addr(Cache_1_io_out_coh_req_bits_addr),
    .io_out_coh_req_bits_wdata(Cache_1_io_out_coh_req_bits_wdata),
    .io_out_coh_resp_valid(Cache_1_io_out_coh_resp_valid),
    .io_out_coh_resp_bits_cmd(Cache_1_io_out_coh_resp_bits_cmd),
    .io_out_coh_resp_bits_rdata(Cache_1_io_out_coh_resp_bits_rdata),
    .io_mmio_req_ready(Cache_1_io_mmio_req_ready),
    .io_mmio_req_valid(Cache_1_io_mmio_req_valid),
    .io_mmio_req_bits_addr(Cache_1_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size(Cache_1_io_mmio_req_bits_size),
    .io_mmio_req_bits_cmd(Cache_1_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(Cache_1_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(Cache_1_io_mmio_req_bits_wdata),
    .io_mmio_resp_valid(Cache_1_io_mmio_resp_valid),
    .io_mmio_resp_bits_rdata(Cache_1_io_mmio_resp_bits_rdata)
  );
  assign io_imem_mem_req_valid = Cache_io_out_mem_req_valid; // @[NutCore.scala 153:13]
  assign io_imem_mem_req_bits_addr = Cache_io_out_mem_req_bits_addr; // @[NutCore.scala 153:13]
  assign io_imem_mem_req_bits_cmd = Cache_io_out_mem_req_bits_cmd; // @[NutCore.scala 153:13]
  assign io_imem_mem_req_bits_wdata = Cache_io_out_mem_req_bits_wdata; // @[NutCore.scala 153:13]
  assign io_dmem_mem_req_valid = Cache_1_io_out_mem_req_valid; // @[NutCore.scala 158:13]
  assign io_dmem_mem_req_bits_addr = Cache_1_io_out_mem_req_bits_addr; // @[NutCore.scala 158:13]
  assign io_dmem_mem_req_bits_cmd = Cache_1_io_out_mem_req_bits_cmd; // @[NutCore.scala 158:13]
  assign io_dmem_mem_req_bits_wdata = Cache_1_io_out_mem_req_bits_wdata; // @[NutCore.scala 158:13]
  assign io_dmem_coh_req_ready = Cache_1_io_out_coh_req_ready; // @[NutCore.scala 158:13]
  assign io_dmem_coh_resp_valid = Cache_1_io_out_coh_resp_valid; // @[NutCore.scala 158:13]
  assign io_dmem_coh_resp_bits_cmd = Cache_1_io_out_coh_resp_bits_cmd; // @[NutCore.scala 158:13]
  assign io_dmem_coh_resp_bits_rdata = Cache_1_io_out_coh_resp_bits_rdata; // @[NutCore.scala 158:13]
  assign io_mmio_req_valid = SimpleBusCrossbarNto1_io_out_req_valid; // @[NutCore.scala 167:13]
  assign io_mmio_req_bits_addr = SimpleBusCrossbarNto1_io_out_req_bits_addr; // @[NutCore.scala 167:13]
  assign io_mmio_req_bits_size = SimpleBusCrossbarNto1_io_out_req_bits_size; // @[NutCore.scala 167:13]
  assign io_mmio_req_bits_cmd = SimpleBusCrossbarNto1_io_out_req_bits_cmd; // @[NutCore.scala 167:13]
  assign io_mmio_req_bits_wmask = SimpleBusCrossbarNto1_io_out_req_bits_wmask; // @[NutCore.scala 167:13]
  assign io_mmio_req_bits_wdata = SimpleBusCrossbarNto1_io_out_req_bits_wdata; // @[NutCore.scala 167:13]
  assign io_frontend_req_ready = SimpleBusCrossbarNto1_1_io_in_3_req_ready; // @[NutCore.scala 165:23]
  assign io_frontend_resp_valid = SimpleBusCrossbarNto1_1_io_in_3_resp_valid; // @[NutCore.scala 165:23]
  assign io_frontend_resp_bits_cmd = SimpleBusCrossbarNto1_1_io_in_3_resp_bits_cmd; // @[NutCore.scala 165:23]
  assign io_frontend_resp_bits_rdata = SimpleBusCrossbarNto1_1_io_in_3_resp_bits_rdata; // @[NutCore.scala 165:23]
  assign perfCnts_2 = Backend_inorder_perfCnts_2;
  assign io_in_bits_decode_cf_pc = Backend_inorder_io_in_bits_decode_cf_pc;
  assign io_wb_rfDest = Backend_inorder_io_wb_rfDest;
  assign io_wb_rfWen = Backend_inorder_io_wb_rfWen;
  assign io_wb_rfData = Backend_inorder_io_wb_rfData;
  assign io_in_valid_0 = Backend_inorder_io_in_valid_0;
  assign frontend_clock = clock;
  assign frontend_reset = reset;
  assign frontend_io_out_0_ready = _T_17 | _T_32; // @[PipelineVector.scala 50:15]
  assign frontend_io_imem_req_ready = EmbeddedTLB_io_in_req_ready; // @[EmbeddedTLB.scala 428:17]
  assign frontend_io_imem_resp_valid = EmbeddedTLB_io_in_resp_valid; // @[EmbeddedTLB.scala 428:17]
  assign frontend_io_imem_resp_bits_rdata = EmbeddedTLB_io_in_resp_bits_rdata; // @[EmbeddedTLB.scala 428:17]
  assign frontend_io_imem_resp_bits_user = EmbeddedTLB_io_in_resp_bits_user; // @[EmbeddedTLB.scala 428:17]
  assign frontend_io_ipf = EmbeddedTLB_io_ipf; // @[NutCore.scala 152:21]
  assign frontend_io_redirect_target = Backend_inorder_io_redirect_target; // @[NutCore.scala 161:26]
  assign frontend_io_redirect_valid = Backend_inorder_io_redirect_valid; // @[NutCore.scala 161:26]
  assign frontend_flushICache = Backend_inorder_flushICache;
  assign frontend__T_243_valid = Backend_inorder__T_243_valid;
  assign frontend__T_243_pc = Backend_inorder__T_243_pc;
  assign frontend__T_243_isMissPredict = Backend_inorder__T_243_isMissPredict;
  assign frontend__T_243_actualTarget = Backend_inorder__T_243_actualTarget;
  assign frontend__T_243_actualTaken = Backend_inorder__T_243_actualTaken;
  assign frontend__T_243_fuOpType = Backend_inorder__T_243_fuOpType;
  assign frontend__T_243_btbType = Backend_inorder__T_243_btbType;
  assign frontend__T_243_isRVC = Backend_inorder__T_243_isRVC;
  assign frontend_vmEnable = EmbeddedTLB_1_vmEnable_0;
  assign frontend_intrVec = Backend_inorder_intrVec;
  assign frontend_flushTLB = Backend_inorder_flushTLB;
  assign Backend_inorder_clock = clock;
  assign Backend_inorder_reset = reset;
  assign Backend_inorder_io_in_0_valid = _T_7 != _T_8; // @[PipelineVector.scala 56:16]
  assign Backend_inorder_io_in_0_bits_cf_instr = 2'h3 == _T_8 ? _T_6_3_cf_instr : _GEN_1167; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_pc = 2'h3 == _T_8 ? _T_6_3_cf_pc : _GEN_1168; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_pnpc = 2'h3 == _T_8 ? _T_6_3_cf_pnpc : _GEN_1169; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_exceptionVec_1 = 2'h3 == _T_8 ? _T_6_3_cf_exceptionVec_1 : _GEN_1174; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_exceptionVec_2 = 2'h3 == _T_8 ? _T_6_3_cf_exceptionVec_2 : _GEN_1175; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_exceptionVec_12 = 2'h3 == _T_8 ? _T_6_3_cf_exceptionVec_12 : _GEN_1185; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_0 = 2'h3 == _T_8 ? _T_6_3_cf_intrVec_0 : _GEN_1189; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_1 = 2'h3 == _T_8 ? _T_6_3_cf_intrVec_1 : _GEN_1190; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_2 = 2'h3 == _T_8 ? _T_6_3_cf_intrVec_2 : _GEN_1191; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_3 = 2'h3 == _T_8 ? _T_6_3_cf_intrVec_3 : _GEN_1192; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_4 = 2'h3 == _T_8 ? _T_6_3_cf_intrVec_4 : _GEN_1193; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_5 = 2'h3 == _T_8 ? _T_6_3_cf_intrVec_5 : _GEN_1194; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_6 = 2'h3 == _T_8 ? _T_6_3_cf_intrVec_6 : _GEN_1195; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_7 = 2'h3 == _T_8 ? _T_6_3_cf_intrVec_7 : _GEN_1196; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_8 = 2'h3 == _T_8 ? _T_6_3_cf_intrVec_8 : _GEN_1197; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_9 = 2'h3 == _T_8 ? _T_6_3_cf_intrVec_9 : _GEN_1198; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_10 = 2'h3 == _T_8 ? _T_6_3_cf_intrVec_10 : _GEN_1199; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_intrVec_11 = 2'h3 == _T_8 ? _T_6_3_cf_intrVec_11 : _GEN_1200; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_brIdx = 2'h3 == _T_8 ? _T_6_3_cf_brIdx : _GEN_1201; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_cf_crossPageIPFFix = 2'h3 == _T_8 ? _T_6_3_cf_crossPageIPFFix : _GEN_1203; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_ctrl_src1Type = 2'h3 == _T_8 ? _T_6_3_ctrl_src1Type : _GEN_1204; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_ctrl_src2Type = 2'h3 == _T_8 ? _T_6_3_ctrl_src2Type : _GEN_1205; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_ctrl_fuType = 2'h3 == _T_8 ? _T_6_3_ctrl_fuType : _GEN_1206; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_ctrl_fuOpType = 2'h3 == _T_8 ? _T_6_3_ctrl_fuOpType : _GEN_1207; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_ctrl_rfSrc1 = 2'h3 == _T_8 ? _T_6_3_ctrl_rfSrc1 : _GEN_1208; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_ctrl_rfSrc2 = 2'h3 == _T_8 ? _T_6_3_ctrl_rfSrc2 : _GEN_1209; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_ctrl_rfWen = 2'h3 == _T_8 ? _T_6_3_ctrl_rfWen : _GEN_1210; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_ctrl_rfDest = 2'h3 == _T_8 ? _T_6_3_ctrl_rfDest : _GEN_1211; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_in_0_bits_data_imm = 2'h3 == _T_8 ? _T_6_3_data_imm : _GEN_1219; // @[PipelineVector.scala 55:15]
  assign Backend_inorder_io_flush = frontend_io_flushVec[3:2]; // @[NutCore.scala 162:22]
  assign Backend_inorder_io_dmem_req_ready = EmbeddedTLB_1_io_in_req_ready; // @[EmbeddedTLB.scala 428:17]
  assign Backend_inorder_io_dmem_resp_valid = EmbeddedTLB_1_io_in_resp_valid; // @[EmbeddedTLB.scala 428:17]
  assign Backend_inorder_io_dmem_resp_bits_rdata = EmbeddedTLB_1_io_in_resp_bits_rdata; // @[EmbeddedTLB.scala 428:17]
  assign Backend_inorder_io_memMMU_dmem_loadPF = EmbeddedTLB_1_io_csrMMU_loadPF; // @[EmbeddedTLB.scala 431:21]
  assign Backend_inorder_io_memMMU_dmem_storePF = EmbeddedTLB_1_io_csrMMU_storePF; // @[EmbeddedTLB.scala 431:21]
  assign Backend_inorder_io_memMMU_dmem_addr = EmbeddedTLB_1_io_csrMMU_addr; // @[EmbeddedTLB.scala 431:21]
  assign Backend_inorder__T_38 = EmbeddedTLB_1__T_38_0;
  assign Backend_inorder_io_extra_mtip = io_extra_mtip;
  assign Backend_inorder_io_extra_meip_0 = io_extra_meip_0;
  assign Backend_inorder_vmEnable = EmbeddedTLB_1_vmEnable_0;
  assign Backend_inorder__T_37 = EmbeddedTLB_1__T_37_0;
  assign Backend_inorder_io_extra_msip = io_extra_msip;
  assign SimpleBusCrossbarNto1_clock = clock;
  assign SimpleBusCrossbarNto1_reset = reset;
  assign SimpleBusCrossbarNto1_io_in_0_req_valid = Cache_io_mmio_req_valid; // @[Cache.scala 685:13]
  assign SimpleBusCrossbarNto1_io_in_0_req_bits_addr = Cache_io_mmio_req_bits_addr; // @[Cache.scala 685:13]
  assign SimpleBusCrossbarNto1_io_in_0_req_bits_cmd = 4'h0; // @[Cache.scala 685:13]
  assign SimpleBusCrossbarNto1_io_in_0_req_bits_wmask = 8'h0; // @[Cache.scala 685:13]
  assign SimpleBusCrossbarNto1_io_in_0_req_bits_wdata = 64'h0; // @[Cache.scala 685:13]
  assign SimpleBusCrossbarNto1_io_in_1_req_valid = Cache_1_io_mmio_req_valid; // @[Cache.scala 685:13]
  assign SimpleBusCrossbarNto1_io_in_1_req_bits_addr = Cache_1_io_mmio_req_bits_addr; // @[Cache.scala 685:13]
  assign SimpleBusCrossbarNto1_io_in_1_req_bits_size = Cache_1_io_mmio_req_bits_size; // @[Cache.scala 685:13]
  assign SimpleBusCrossbarNto1_io_in_1_req_bits_cmd = Cache_1_io_mmio_req_bits_cmd; // @[Cache.scala 685:13]
  assign SimpleBusCrossbarNto1_io_in_1_req_bits_wmask = Cache_1_io_mmio_req_bits_wmask; // @[Cache.scala 685:13]
  assign SimpleBusCrossbarNto1_io_in_1_req_bits_wdata = Cache_1_io_mmio_req_bits_wdata; // @[Cache.scala 685:13]
  assign SimpleBusCrossbarNto1_io_out_req_ready = io_mmio_req_ready; // @[NutCore.scala 167:13]
  assign SimpleBusCrossbarNto1_io_out_resp_valid = io_mmio_resp_valid; // @[NutCore.scala 167:13]
  assign SimpleBusCrossbarNto1_io_out_resp_bits_cmd = io_mmio_resp_bits_cmd; // @[NutCore.scala 167:13]
  assign SimpleBusCrossbarNto1_io_out_resp_bits_rdata = io_mmio_resp_bits_rdata; // @[NutCore.scala 167:13]
  assign SimpleBusCrossbarNto1_1_clock = clock;
  assign SimpleBusCrossbarNto1_1_reset = reset;
  assign SimpleBusCrossbarNto1_1_io_in_0_req_valid = EmbeddedTLB_1_io_out_req_valid; // @[NutCore.scala 157:23]
  assign SimpleBusCrossbarNto1_1_io_in_0_req_bits_addr = EmbeddedTLB_1_io_out_req_bits_addr; // @[NutCore.scala 157:23]
  assign SimpleBusCrossbarNto1_1_io_in_0_req_bits_size = EmbeddedTLB_1_io_out_req_bits_size; // @[NutCore.scala 157:23]
  assign SimpleBusCrossbarNto1_1_io_in_0_req_bits_cmd = EmbeddedTLB_1_io_out_req_bits_cmd; // @[NutCore.scala 157:23]
  assign SimpleBusCrossbarNto1_1_io_in_0_req_bits_wmask = EmbeddedTLB_1_io_out_req_bits_wmask; // @[NutCore.scala 157:23]
  assign SimpleBusCrossbarNto1_1_io_in_0_req_bits_wdata = EmbeddedTLB_1_io_out_req_bits_wdata; // @[NutCore.scala 157:23]
  assign SimpleBusCrossbarNto1_1_io_in_1_req_valid = EmbeddedTLB_io_mem_req_valid; // @[EmbeddedTLB.scala 429:18]
  assign SimpleBusCrossbarNto1_1_io_in_1_req_bits_addr = EmbeddedTLB_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 429:18]
  assign SimpleBusCrossbarNto1_1_io_in_1_req_bits_cmd = EmbeddedTLB_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 429:18]
  assign SimpleBusCrossbarNto1_1_io_in_1_req_bits_wdata = EmbeddedTLB_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 429:18]
  assign SimpleBusCrossbarNto1_1_io_in_2_req_valid = EmbeddedTLB_1_io_mem_req_valid; // @[EmbeddedTLB.scala 429:18]
  assign SimpleBusCrossbarNto1_1_io_in_2_req_bits_addr = EmbeddedTLB_1_io_mem_req_bits_addr; // @[EmbeddedTLB.scala 429:18]
  assign SimpleBusCrossbarNto1_1_io_in_2_req_bits_cmd = EmbeddedTLB_1_io_mem_req_bits_cmd; // @[EmbeddedTLB.scala 429:18]
  assign SimpleBusCrossbarNto1_1_io_in_2_req_bits_wdata = EmbeddedTLB_1_io_mem_req_bits_wdata; // @[EmbeddedTLB.scala 429:18]
  assign SimpleBusCrossbarNto1_1_io_in_3_req_valid = io_frontend_req_valid; // @[NutCore.scala 165:23]
  assign SimpleBusCrossbarNto1_1_io_in_3_req_bits_addr = io_frontend_req_bits_addr; // @[NutCore.scala 165:23]
  assign SimpleBusCrossbarNto1_1_io_in_3_req_bits_size = io_frontend_req_bits_size; // @[NutCore.scala 165:23]
  assign SimpleBusCrossbarNto1_1_io_in_3_req_bits_cmd = io_frontend_req_bits_cmd; // @[NutCore.scala 165:23]
  assign SimpleBusCrossbarNto1_1_io_in_3_req_bits_wmask = io_frontend_req_bits_wmask; // @[NutCore.scala 165:23]
  assign SimpleBusCrossbarNto1_1_io_in_3_req_bits_wdata = io_frontend_req_bits_wdata; // @[NutCore.scala 165:23]
  assign SimpleBusCrossbarNto1_1_io_in_3_resp_ready = io_frontend_resp_ready; // @[NutCore.scala 165:23]
  assign SimpleBusCrossbarNto1_1_io_out_req_ready = Cache_1_io_in_req_ready; // @[Cache.scala 684:17]
  assign SimpleBusCrossbarNto1_1_io_out_resp_valid = Cache_1_io_in_resp_valid; // @[Cache.scala 684:17]
  assign SimpleBusCrossbarNto1_1_io_out_resp_bits_cmd = Cache_1_io_in_resp_bits_cmd; // @[Cache.scala 684:17]
  assign SimpleBusCrossbarNto1_1_io_out_resp_bits_rdata = Cache_1_io_in_resp_bits_rdata; // @[Cache.scala 684:17]
  assign EmbeddedTLB_clock = clock;
  assign EmbeddedTLB_reset = reset;
  assign EmbeddedTLB_io_in_req_valid = frontend_io_imem_req_valid; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_io_in_req_bits_addr = frontend_io_imem_req_bits_addr; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_io_in_req_bits_user = frontend_io_imem_req_bits_user; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_io_in_resp_ready = frontend_io_imem_resp_ready; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_io_out_req_ready = Cache_io_in_req_ready; // @[Cache.scala 684:17]
  assign EmbeddedTLB_io_out_resp_valid = Cache_io_in_resp_valid; // @[Cache.scala 684:17]
  assign EmbeddedTLB_io_out_resp_bits_rdata = Cache_io_in_resp_bits_rdata; // @[Cache.scala 684:17]
  assign EmbeddedTLB_io_out_resp_bits_user = Cache_io_in_resp_bits_user; // @[Cache.scala 684:17]
  assign EmbeddedTLB_io_mem_req_ready = SimpleBusCrossbarNto1_1_io_in_1_req_ready; // @[EmbeddedTLB.scala 429:18]
  assign EmbeddedTLB_io_mem_resp_valid = SimpleBusCrossbarNto1_1_io_in_1_resp_valid; // @[EmbeddedTLB.scala 429:18]
  assign EmbeddedTLB_io_mem_resp_bits_rdata = SimpleBusCrossbarNto1_1_io_in_1_resp_bits_rdata; // @[EmbeddedTLB.scala 429:18]
  assign EmbeddedTLB_io_flush = frontend_io_flushVec[0]; // @[EmbeddedTLB.scala 430:20]
  assign EmbeddedTLB_io_csrMMU_priviledgeMode = Backend_inorder_io_memMMU_imem_priviledgeMode; // @[EmbeddedTLB.scala 431:21]
  assign EmbeddedTLB_io_cacheEmpty = Cache_io_empty; // @[Cache.scala 686:11]
  assign EmbeddedTLB_CSRSATP = Backend_inorder_satp;
  assign EmbeddedTLB_MOUFlushTLB = Backend_inorder_flushTLB;
  assign Cache_clock = clock;
  assign Cache_reset = reset;
  assign Cache_io_in_req_valid = EmbeddedTLB_io_out_req_valid; // @[Cache.scala 684:17]
  assign Cache_io_in_req_bits_addr = EmbeddedTLB_io_out_req_bits_addr; // @[Cache.scala 684:17]
  assign Cache_io_in_req_bits_user = EmbeddedTLB_io_out_req_bits_user; // @[Cache.scala 684:17]
  assign Cache_io_in_resp_ready = EmbeddedTLB_io_out_resp_ready; // @[Cache.scala 684:17]
  assign Cache_io_flush = frontend_io_flushVec[0] ? 2'h3 : 2'h0; // @[Cache.scala 683:20]
  assign Cache_io_out_mem_req_ready = io_imem_mem_req_ready; // @[NutCore.scala 153:13]
  assign Cache_io_out_mem_resp_valid = io_imem_mem_resp_valid; // @[NutCore.scala 153:13]
  assign Cache_io_out_mem_resp_bits_cmd = io_imem_mem_resp_bits_cmd; // @[NutCore.scala 153:13]
  assign Cache_io_out_mem_resp_bits_rdata = io_imem_mem_resp_bits_rdata; // @[NutCore.scala 153:13]
  assign Cache_io_mmio_req_ready = SimpleBusCrossbarNto1_io_in_0_req_ready; // @[Cache.scala 685:13]
  assign Cache_io_mmio_resp_valid = SimpleBusCrossbarNto1_io_in_0_resp_valid; // @[Cache.scala 685:13]
  assign Cache_io_mmio_resp_bits_rdata = SimpleBusCrossbarNto1_io_in_0_resp_bits_rdata; // @[Cache.scala 685:13]
  assign Cache_MOUFlushICache = Backend_inorder_flushICache;
  assign EmbeddedTLB_1_clock = clock;
  assign EmbeddedTLB_1_reset = reset;
  assign EmbeddedTLB_1_io_in_req_valid = Backend_inorder_io_dmem_req_valid; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_1_io_in_req_bits_addr = Backend_inorder_io_dmem_req_bits_addr; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_1_io_in_req_bits_size = Backend_inorder_io_dmem_req_bits_size; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_1_io_in_req_bits_cmd = Backend_inorder_io_dmem_req_bits_cmd; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_1_io_in_req_bits_wmask = Backend_inorder_io_dmem_req_bits_wmask; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_1_io_in_req_bits_wdata = Backend_inorder_io_dmem_req_bits_wdata; // @[EmbeddedTLB.scala 428:17]
  assign EmbeddedTLB_1_io_out_req_ready = SimpleBusCrossbarNto1_1_io_in_0_req_ready; // @[NutCore.scala 157:23]
  assign EmbeddedTLB_1_io_out_resp_valid = SimpleBusCrossbarNto1_1_io_in_0_resp_valid; // @[NutCore.scala 157:23]
  assign EmbeddedTLB_1_io_out_resp_bits_rdata = SimpleBusCrossbarNto1_1_io_in_0_resp_bits_rdata; // @[NutCore.scala 157:23]
  assign EmbeddedTLB_1_io_mem_req_ready = SimpleBusCrossbarNto1_1_io_in_2_req_ready; // @[EmbeddedTLB.scala 429:18]
  assign EmbeddedTLB_1_io_mem_resp_valid = SimpleBusCrossbarNto1_1_io_in_2_resp_valid; // @[EmbeddedTLB.scala 429:18]
  assign EmbeddedTLB_1_io_mem_resp_bits_rdata = SimpleBusCrossbarNto1_1_io_in_2_resp_bits_rdata; // @[EmbeddedTLB.scala 429:18]
  assign EmbeddedTLB_1_io_csrMMU_priviledgeMode = Backend_inorder_io_memMMU_dmem_priviledgeMode; // @[EmbeddedTLB.scala 431:21]
  assign EmbeddedTLB_1_io_csrMMU_status_sum = Backend_inorder_io_memMMU_dmem_status_sum; // @[EmbeddedTLB.scala 431:21]
  assign EmbeddedTLB_1_io_csrMMU_status_mxr = Backend_inorder_io_memMMU_dmem_status_mxr; // @[EmbeddedTLB.scala 431:21]
  assign EmbeddedTLB_1_CSRSATP = Backend_inorder_satp;
  assign EmbeddedTLB_1_amoReq = Backend_inorder_amoReq;
  assign EmbeddedTLB_1_MOUFlushTLB = Backend_inorder_flushTLB;
  assign Cache_1_clock = clock;
  assign Cache_1_reset = reset;
  assign Cache_1_io_in_req_valid = SimpleBusCrossbarNto1_1_io_out_req_valid; // @[Cache.scala 684:17]
  assign Cache_1_io_in_req_bits_addr = SimpleBusCrossbarNto1_1_io_out_req_bits_addr; // @[Cache.scala 684:17]
  assign Cache_1_io_in_req_bits_size = SimpleBusCrossbarNto1_1_io_out_req_bits_size; // @[Cache.scala 684:17]
  assign Cache_1_io_in_req_bits_cmd = SimpleBusCrossbarNto1_1_io_out_req_bits_cmd; // @[Cache.scala 684:17]
  assign Cache_1_io_in_req_bits_wmask = SimpleBusCrossbarNto1_1_io_out_req_bits_wmask; // @[Cache.scala 684:17]
  assign Cache_1_io_in_req_bits_wdata = SimpleBusCrossbarNto1_1_io_out_req_bits_wdata; // @[Cache.scala 684:17]
  assign Cache_1_io_in_resp_ready = SimpleBusCrossbarNto1_1_io_out_resp_ready; // @[Cache.scala 684:17]
  assign Cache_1_io_out_mem_req_ready = io_dmem_mem_req_ready; // @[NutCore.scala 158:13]
  assign Cache_1_io_out_mem_resp_valid = io_dmem_mem_resp_valid; // @[NutCore.scala 158:13]
  assign Cache_1_io_out_mem_resp_bits_cmd = io_dmem_mem_resp_bits_cmd; // @[NutCore.scala 158:13]
  assign Cache_1_io_out_mem_resp_bits_rdata = io_dmem_mem_resp_bits_rdata; // @[NutCore.scala 158:13]
  assign Cache_1_io_out_coh_req_valid = io_dmem_coh_req_valid; // @[NutCore.scala 158:13]
  assign Cache_1_io_out_coh_req_bits_addr = io_dmem_coh_req_bits_addr; // @[NutCore.scala 158:13]
  assign Cache_1_io_out_coh_req_bits_wdata = io_dmem_coh_req_bits_wdata; // @[NutCore.scala 158:13]
  assign Cache_1_io_mmio_req_ready = SimpleBusCrossbarNto1_io_in_1_req_ready; // @[Cache.scala 685:13]
  assign Cache_1_io_mmio_resp_valid = SimpleBusCrossbarNto1_io_in_1_resp_valid; // @[Cache.scala 685:13]
  assign Cache_1_io_mmio_resp_bits_rdata = SimpleBusCrossbarNto1_io_in_1_resp_bits_rdata; // @[Cache.scala 685:13]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {2{`RANDOM}};
  _T_6_0_cf_instr = _RAND_0[63:0];
  _RAND_1 = {2{`RANDOM}};
  _T_6_0_cf_pc = _RAND_1[38:0];
  _RAND_2 = {2{`RANDOM}};
  _T_6_0_cf_pnpc = _RAND_2[38:0];
  _RAND_3 = {1{`RANDOM}};
  _T_6_0_cf_exceptionVec_1 = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_6_0_cf_exceptionVec_2 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  _T_6_0_cf_exceptionVec_12 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_6_0_cf_intrVec_0 = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_6_0_cf_intrVec_1 = _RAND_7[0:0];
  _RAND_8 = {1{`RANDOM}};
  _T_6_0_cf_intrVec_2 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _T_6_0_cf_intrVec_3 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _T_6_0_cf_intrVec_4 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  _T_6_0_cf_intrVec_5 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _T_6_0_cf_intrVec_6 = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _T_6_0_cf_intrVec_7 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  _T_6_0_cf_intrVec_8 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _T_6_0_cf_intrVec_9 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  _T_6_0_cf_intrVec_10 = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  _T_6_0_cf_intrVec_11 = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _T_6_0_cf_brIdx = _RAND_18[3:0];
  _RAND_19 = {1{`RANDOM}};
  _T_6_0_cf_crossPageIPFFix = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  _T_6_0_ctrl_src1Type = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _T_6_0_ctrl_src2Type = _RAND_21[0:0];
  _RAND_22 = {1{`RANDOM}};
  _T_6_0_ctrl_fuType = _RAND_22[2:0];
  _RAND_23 = {1{`RANDOM}};
  _T_6_0_ctrl_fuOpType = _RAND_23[6:0];
  _RAND_24 = {1{`RANDOM}};
  _T_6_0_ctrl_rfSrc1 = _RAND_24[4:0];
  _RAND_25 = {1{`RANDOM}};
  _T_6_0_ctrl_rfSrc2 = _RAND_25[4:0];
  _RAND_26 = {1{`RANDOM}};
  _T_6_0_ctrl_rfWen = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  _T_6_0_ctrl_rfDest = _RAND_27[4:0];
  _RAND_28 = {2{`RANDOM}};
  _T_6_0_data_imm = _RAND_28[63:0];
  _RAND_29 = {2{`RANDOM}};
  _T_6_1_cf_instr = _RAND_29[63:0];
  _RAND_30 = {2{`RANDOM}};
  _T_6_1_cf_pc = _RAND_30[38:0];
  _RAND_31 = {2{`RANDOM}};
  _T_6_1_cf_pnpc = _RAND_31[38:0];
  _RAND_32 = {1{`RANDOM}};
  _T_6_1_cf_exceptionVec_1 = _RAND_32[0:0];
  _RAND_33 = {1{`RANDOM}};
  _T_6_1_cf_exceptionVec_2 = _RAND_33[0:0];
  _RAND_34 = {1{`RANDOM}};
  _T_6_1_cf_exceptionVec_12 = _RAND_34[0:0];
  _RAND_35 = {1{`RANDOM}};
  _T_6_1_cf_intrVec_0 = _RAND_35[0:0];
  _RAND_36 = {1{`RANDOM}};
  _T_6_1_cf_intrVec_1 = _RAND_36[0:0];
  _RAND_37 = {1{`RANDOM}};
  _T_6_1_cf_intrVec_2 = _RAND_37[0:0];
  _RAND_38 = {1{`RANDOM}};
  _T_6_1_cf_intrVec_3 = _RAND_38[0:0];
  _RAND_39 = {1{`RANDOM}};
  _T_6_1_cf_intrVec_4 = _RAND_39[0:0];
  _RAND_40 = {1{`RANDOM}};
  _T_6_1_cf_intrVec_5 = _RAND_40[0:0];
  _RAND_41 = {1{`RANDOM}};
  _T_6_1_cf_intrVec_6 = _RAND_41[0:0];
  _RAND_42 = {1{`RANDOM}};
  _T_6_1_cf_intrVec_7 = _RAND_42[0:0];
  _RAND_43 = {1{`RANDOM}};
  _T_6_1_cf_intrVec_8 = _RAND_43[0:0];
  _RAND_44 = {1{`RANDOM}};
  _T_6_1_cf_intrVec_9 = _RAND_44[0:0];
  _RAND_45 = {1{`RANDOM}};
  _T_6_1_cf_intrVec_10 = _RAND_45[0:0];
  _RAND_46 = {1{`RANDOM}};
  _T_6_1_cf_intrVec_11 = _RAND_46[0:0];
  _RAND_47 = {1{`RANDOM}};
  _T_6_1_cf_brIdx = _RAND_47[3:0];
  _RAND_48 = {1{`RANDOM}};
  _T_6_1_cf_crossPageIPFFix = _RAND_48[0:0];
  _RAND_49 = {1{`RANDOM}};
  _T_6_1_ctrl_src1Type = _RAND_49[0:0];
  _RAND_50 = {1{`RANDOM}};
  _T_6_1_ctrl_src2Type = _RAND_50[0:0];
  _RAND_51 = {1{`RANDOM}};
  _T_6_1_ctrl_fuType = _RAND_51[2:0];
  _RAND_52 = {1{`RANDOM}};
  _T_6_1_ctrl_fuOpType = _RAND_52[6:0];
  _RAND_53 = {1{`RANDOM}};
  _T_6_1_ctrl_rfSrc1 = _RAND_53[4:0];
  _RAND_54 = {1{`RANDOM}};
  _T_6_1_ctrl_rfSrc2 = _RAND_54[4:0];
  _RAND_55 = {1{`RANDOM}};
  _T_6_1_ctrl_rfWen = _RAND_55[0:0];
  _RAND_56 = {1{`RANDOM}};
  _T_6_1_ctrl_rfDest = _RAND_56[4:0];
  _RAND_57 = {2{`RANDOM}};
  _T_6_1_data_imm = _RAND_57[63:0];
  _RAND_58 = {2{`RANDOM}};
  _T_6_2_cf_instr = _RAND_58[63:0];
  _RAND_59 = {2{`RANDOM}};
  _T_6_2_cf_pc = _RAND_59[38:0];
  _RAND_60 = {2{`RANDOM}};
  _T_6_2_cf_pnpc = _RAND_60[38:0];
  _RAND_61 = {1{`RANDOM}};
  _T_6_2_cf_exceptionVec_1 = _RAND_61[0:0];
  _RAND_62 = {1{`RANDOM}};
  _T_6_2_cf_exceptionVec_2 = _RAND_62[0:0];
  _RAND_63 = {1{`RANDOM}};
  _T_6_2_cf_exceptionVec_12 = _RAND_63[0:0];
  _RAND_64 = {1{`RANDOM}};
  _T_6_2_cf_intrVec_0 = _RAND_64[0:0];
  _RAND_65 = {1{`RANDOM}};
  _T_6_2_cf_intrVec_1 = _RAND_65[0:0];
  _RAND_66 = {1{`RANDOM}};
  _T_6_2_cf_intrVec_2 = _RAND_66[0:0];
  _RAND_67 = {1{`RANDOM}};
  _T_6_2_cf_intrVec_3 = _RAND_67[0:0];
  _RAND_68 = {1{`RANDOM}};
  _T_6_2_cf_intrVec_4 = _RAND_68[0:0];
  _RAND_69 = {1{`RANDOM}};
  _T_6_2_cf_intrVec_5 = _RAND_69[0:0];
  _RAND_70 = {1{`RANDOM}};
  _T_6_2_cf_intrVec_6 = _RAND_70[0:0];
  _RAND_71 = {1{`RANDOM}};
  _T_6_2_cf_intrVec_7 = _RAND_71[0:0];
  _RAND_72 = {1{`RANDOM}};
  _T_6_2_cf_intrVec_8 = _RAND_72[0:0];
  _RAND_73 = {1{`RANDOM}};
  _T_6_2_cf_intrVec_9 = _RAND_73[0:0];
  _RAND_74 = {1{`RANDOM}};
  _T_6_2_cf_intrVec_10 = _RAND_74[0:0];
  _RAND_75 = {1{`RANDOM}};
  _T_6_2_cf_intrVec_11 = _RAND_75[0:0];
  _RAND_76 = {1{`RANDOM}};
  _T_6_2_cf_brIdx = _RAND_76[3:0];
  _RAND_77 = {1{`RANDOM}};
  _T_6_2_cf_crossPageIPFFix = _RAND_77[0:0];
  _RAND_78 = {1{`RANDOM}};
  _T_6_2_ctrl_src1Type = _RAND_78[0:0];
  _RAND_79 = {1{`RANDOM}};
  _T_6_2_ctrl_src2Type = _RAND_79[0:0];
  _RAND_80 = {1{`RANDOM}};
  _T_6_2_ctrl_fuType = _RAND_80[2:0];
  _RAND_81 = {1{`RANDOM}};
  _T_6_2_ctrl_fuOpType = _RAND_81[6:0];
  _RAND_82 = {1{`RANDOM}};
  _T_6_2_ctrl_rfSrc1 = _RAND_82[4:0];
  _RAND_83 = {1{`RANDOM}};
  _T_6_2_ctrl_rfSrc2 = _RAND_83[4:0];
  _RAND_84 = {1{`RANDOM}};
  _T_6_2_ctrl_rfWen = _RAND_84[0:0];
  _RAND_85 = {1{`RANDOM}};
  _T_6_2_ctrl_rfDest = _RAND_85[4:0];
  _RAND_86 = {2{`RANDOM}};
  _T_6_2_data_imm = _RAND_86[63:0];
  _RAND_87 = {2{`RANDOM}};
  _T_6_3_cf_instr = _RAND_87[63:0];
  _RAND_88 = {2{`RANDOM}};
  _T_6_3_cf_pc = _RAND_88[38:0];
  _RAND_89 = {2{`RANDOM}};
  _T_6_3_cf_pnpc = _RAND_89[38:0];
  _RAND_90 = {1{`RANDOM}};
  _T_6_3_cf_exceptionVec_1 = _RAND_90[0:0];
  _RAND_91 = {1{`RANDOM}};
  _T_6_3_cf_exceptionVec_2 = _RAND_91[0:0];
  _RAND_92 = {1{`RANDOM}};
  _T_6_3_cf_exceptionVec_12 = _RAND_92[0:0];
  _RAND_93 = {1{`RANDOM}};
  _T_6_3_cf_intrVec_0 = _RAND_93[0:0];
  _RAND_94 = {1{`RANDOM}};
  _T_6_3_cf_intrVec_1 = _RAND_94[0:0];
  _RAND_95 = {1{`RANDOM}};
  _T_6_3_cf_intrVec_2 = _RAND_95[0:0];
  _RAND_96 = {1{`RANDOM}};
  _T_6_3_cf_intrVec_3 = _RAND_96[0:0];
  _RAND_97 = {1{`RANDOM}};
  _T_6_3_cf_intrVec_4 = _RAND_97[0:0];
  _RAND_98 = {1{`RANDOM}};
  _T_6_3_cf_intrVec_5 = _RAND_98[0:0];
  _RAND_99 = {1{`RANDOM}};
  _T_6_3_cf_intrVec_6 = _RAND_99[0:0];
  _RAND_100 = {1{`RANDOM}};
  _T_6_3_cf_intrVec_7 = _RAND_100[0:0];
  _RAND_101 = {1{`RANDOM}};
  _T_6_3_cf_intrVec_8 = _RAND_101[0:0];
  _RAND_102 = {1{`RANDOM}};
  _T_6_3_cf_intrVec_9 = _RAND_102[0:0];
  _RAND_103 = {1{`RANDOM}};
  _T_6_3_cf_intrVec_10 = _RAND_103[0:0];
  _RAND_104 = {1{`RANDOM}};
  _T_6_3_cf_intrVec_11 = _RAND_104[0:0];
  _RAND_105 = {1{`RANDOM}};
  _T_6_3_cf_brIdx = _RAND_105[3:0];
  _RAND_106 = {1{`RANDOM}};
  _T_6_3_cf_crossPageIPFFix = _RAND_106[0:0];
  _RAND_107 = {1{`RANDOM}};
  _T_6_3_ctrl_src1Type = _RAND_107[0:0];
  _RAND_108 = {1{`RANDOM}};
  _T_6_3_ctrl_src2Type = _RAND_108[0:0];
  _RAND_109 = {1{`RANDOM}};
  _T_6_3_ctrl_fuType = _RAND_109[2:0];
  _RAND_110 = {1{`RANDOM}};
  _T_6_3_ctrl_fuOpType = _RAND_110[6:0];
  _RAND_111 = {1{`RANDOM}};
  _T_6_3_ctrl_rfSrc1 = _RAND_111[4:0];
  _RAND_112 = {1{`RANDOM}};
  _T_6_3_ctrl_rfSrc2 = _RAND_112[4:0];
  _RAND_113 = {1{`RANDOM}};
  _T_6_3_ctrl_rfWen = _RAND_113[0:0];
  _RAND_114 = {1{`RANDOM}};
  _T_6_3_ctrl_rfDest = _RAND_114[4:0];
  _RAND_115 = {2{`RANDOM}};
  _T_6_3_data_imm = _RAND_115[63:0];
  _RAND_116 = {1{`RANDOM}};
  _T_7 = _RAND_116[1:0];
  _RAND_117 = {1{`RANDOM}};
  _T_8 = _RAND_117[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_6_0_cf_instr <= 64'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_instr <= 64'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_instr <= frontend_io_out_0_bits_cf_instr;
            end else begin
              _T_6_0_cf_instr <= 64'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_instr <= frontend_io_out_0_bits_cf_instr;
          end else begin
            _T_6_0_cf_instr <= 64'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_pc <= 39'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_pc <= 39'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_pc <= frontend_io_out_0_bits_cf_pc;
            end else begin
              _T_6_0_cf_pc <= 39'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_pc <= frontend_io_out_0_bits_cf_pc;
          end else begin
            _T_6_0_cf_pc <= 39'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_pnpc <= 39'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_pnpc <= 39'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_pnpc <= frontend_io_out_0_bits_cf_pnpc;
            end else begin
              _T_6_0_cf_pnpc <= 39'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_pnpc <= frontend_io_out_0_bits_cf_pnpc;
          end else begin
            _T_6_0_cf_pnpc <= 39'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_exceptionVec_1 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_exceptionVec_1 <= 1'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            _T_6_0_cf_exceptionVec_1 <= _T_27_cf_exceptionVec_1;
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          _T_6_0_cf_exceptionVec_1 <= _T_27_cf_exceptionVec_1;
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_exceptionVec_2 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_exceptionVec_2 <= 1'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            _T_6_0_cf_exceptionVec_2 <= _T_27_cf_exceptionVec_2;
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          _T_6_0_cf_exceptionVec_2 <= _T_27_cf_exceptionVec_2;
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_exceptionVec_12 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_exceptionVec_12 <= 1'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            _T_6_0_cf_exceptionVec_12 <= _T_27_cf_exceptionVec_12;
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          _T_6_0_cf_exceptionVec_12 <= _T_27_cf_exceptionVec_12;
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_intrVec_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_intrVec_0 <= _T_6_T_29_cf_intrVec_0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_intrVec_0 <= frontend_io_out_0_bits_cf_intrVec_0;
            end else begin
              _T_6_0_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_intrVec_0 <= frontend_io_out_0_bits_cf_intrVec_0;
          end else begin
            _T_6_0_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_intrVec_1 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_intrVec_1 <= _T_6_T_29_cf_intrVec_1;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_intrVec_1 <= frontend_io_out_0_bits_cf_intrVec_1;
            end else begin
              _T_6_0_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_intrVec_1 <= frontend_io_out_0_bits_cf_intrVec_1;
          end else begin
            _T_6_0_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_intrVec_2 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_intrVec_2 <= _T_6_T_29_cf_intrVec_2;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_intrVec_2 <= frontend_io_out_0_bits_cf_intrVec_2;
            end else begin
              _T_6_0_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_intrVec_2 <= frontend_io_out_0_bits_cf_intrVec_2;
          end else begin
            _T_6_0_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_intrVec_3 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_intrVec_3 <= _T_6_T_29_cf_intrVec_3;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_intrVec_3 <= frontend_io_out_0_bits_cf_intrVec_3;
            end else begin
              _T_6_0_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_intrVec_3 <= frontend_io_out_0_bits_cf_intrVec_3;
          end else begin
            _T_6_0_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_intrVec_4 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_intrVec_4 <= _T_6_T_29_cf_intrVec_4;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_intrVec_4 <= frontend_io_out_0_bits_cf_intrVec_4;
            end else begin
              _T_6_0_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_intrVec_4 <= frontend_io_out_0_bits_cf_intrVec_4;
          end else begin
            _T_6_0_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_intrVec_5 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_intrVec_5 <= _T_6_T_29_cf_intrVec_5;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_intrVec_5 <= frontend_io_out_0_bits_cf_intrVec_5;
            end else begin
              _T_6_0_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_intrVec_5 <= frontend_io_out_0_bits_cf_intrVec_5;
          end else begin
            _T_6_0_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_intrVec_6 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_intrVec_6 <= _T_6_T_29_cf_intrVec_6;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_intrVec_6 <= frontend_io_out_0_bits_cf_intrVec_6;
            end else begin
              _T_6_0_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_intrVec_6 <= frontend_io_out_0_bits_cf_intrVec_6;
          end else begin
            _T_6_0_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_intrVec_7 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_intrVec_7 <= _T_6_T_29_cf_intrVec_7;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_intrVec_7 <= frontend_io_out_0_bits_cf_intrVec_7;
            end else begin
              _T_6_0_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_intrVec_7 <= frontend_io_out_0_bits_cf_intrVec_7;
          end else begin
            _T_6_0_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_intrVec_8 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_intrVec_8 <= _T_6_T_29_cf_intrVec_8;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_intrVec_8 <= frontend_io_out_0_bits_cf_intrVec_8;
            end else begin
              _T_6_0_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_intrVec_8 <= frontend_io_out_0_bits_cf_intrVec_8;
          end else begin
            _T_6_0_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_intrVec_9 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_intrVec_9 <= _T_6_T_29_cf_intrVec_9;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_intrVec_9 <= frontend_io_out_0_bits_cf_intrVec_9;
            end else begin
              _T_6_0_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_intrVec_9 <= frontend_io_out_0_bits_cf_intrVec_9;
          end else begin
            _T_6_0_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_intrVec_10 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_intrVec_10 <= _T_6_T_29_cf_intrVec_10;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_intrVec_10 <= frontend_io_out_0_bits_cf_intrVec_10;
            end else begin
              _T_6_0_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_intrVec_10 <= frontend_io_out_0_bits_cf_intrVec_10;
          end else begin
            _T_6_0_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_intrVec_11 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_intrVec_11 <= _T_6_T_29_cf_intrVec_11;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_intrVec_11 <= frontend_io_out_0_bits_cf_intrVec_11;
            end else begin
              _T_6_0_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_intrVec_11 <= frontend_io_out_0_bits_cf_intrVec_11;
          end else begin
            _T_6_0_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_brIdx <= 4'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_brIdx <= 4'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_cf_brIdx <= frontend_io_out_0_bits_cf_brIdx;
            end else begin
              _T_6_0_cf_brIdx <= 4'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_cf_brIdx <= frontend_io_out_0_bits_cf_brIdx;
          end else begin
            _T_6_0_cf_brIdx <= 4'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_cf_crossPageIPFFix <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_cf_crossPageIPFFix <= 1'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            _T_6_0_cf_crossPageIPFFix <= _T_27_cf_crossPageIPFFix;
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          _T_6_0_cf_crossPageIPFFix <= _T_27_cf_crossPageIPFFix;
        end
      end
    end
    if (reset) begin
      _T_6_0_ctrl_src1Type <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        _T_6_0_ctrl_src1Type <= _GEN_484;
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_ctrl_src1Type <= frontend_io_out_0_bits_ctrl_src1Type;
          end else begin
            _T_6_0_ctrl_src1Type <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_ctrl_src2Type <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        _T_6_0_ctrl_src2Type <= _GEN_480;
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_ctrl_src2Type <= frontend_io_out_0_bits_ctrl_src2Type;
          end else begin
            _T_6_0_ctrl_src2Type <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_ctrl_fuType <= 3'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_ctrl_fuType <= 3'h3;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_ctrl_fuType <= frontend_io_out_0_bits_ctrl_fuType;
            end else begin
              _T_6_0_ctrl_fuType <= 3'h3;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_ctrl_fuType <= frontend_io_out_0_bits_ctrl_fuType;
          end else begin
            _T_6_0_ctrl_fuType <= 3'h3;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_ctrl_fuOpType <= 7'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_ctrl_fuOpType <= 7'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_ctrl_fuOpType <= frontend_io_out_0_bits_ctrl_fuOpType;
            end else begin
              _T_6_0_ctrl_fuOpType <= 7'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_ctrl_fuOpType <= frontend_io_out_0_bits_ctrl_fuOpType;
          end else begin
            _T_6_0_ctrl_fuOpType <= 7'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_ctrl_rfSrc1 <= 5'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_ctrl_rfSrc1 <= 5'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_ctrl_rfSrc1 <= frontend_io_out_0_bits_ctrl_rfSrc1;
            end else begin
              _T_6_0_ctrl_rfSrc1 <= 5'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_ctrl_rfSrc1 <= frontend_io_out_0_bits_ctrl_rfSrc1;
          end else begin
            _T_6_0_ctrl_rfSrc1 <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_ctrl_rfSrc2 <= 5'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_ctrl_rfSrc2 <= 5'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_ctrl_rfSrc2 <= frontend_io_out_0_bits_ctrl_rfSrc2;
            end else begin
              _T_6_0_ctrl_rfSrc2 <= 5'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_ctrl_rfSrc2 <= frontend_io_out_0_bits_ctrl_rfSrc2;
          end else begin
            _T_6_0_ctrl_rfSrc2 <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_ctrl_rfWen <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_ctrl_rfWen <= 1'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            _T_6_0_ctrl_rfWen <= _T_27_ctrl_rfWen;
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          _T_6_0_ctrl_rfWen <= _T_27_ctrl_rfWen;
        end
      end
    end
    if (reset) begin
      _T_6_0_ctrl_rfDest <= 5'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_ctrl_rfDest <= 5'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_ctrl_rfDest <= frontend_io_out_0_bits_ctrl_rfDest;
            end else begin
              _T_6_0_ctrl_rfDest <= 5'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_ctrl_rfDest <= frontend_io_out_0_bits_ctrl_rfDest;
          end else begin
            _T_6_0_ctrl_rfDest <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_0_data_imm <= 64'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h0 == _T_29) begin
          _T_6_0_data_imm <= 64'h0;
        end else if (_T_20) begin
          if (2'h0 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_0_data_imm <= frontend_io_out_0_bits_data_imm;
            end else begin
              _T_6_0_data_imm <= 64'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h0 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_0_data_imm <= frontend_io_out_0_bits_data_imm;
          end else begin
            _T_6_0_data_imm <= 64'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_instr <= 64'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_instr <= 64'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_instr <= frontend_io_out_0_bits_cf_instr;
            end else begin
              _T_6_1_cf_instr <= 64'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_instr <= frontend_io_out_0_bits_cf_instr;
          end else begin
            _T_6_1_cf_instr <= 64'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_pc <= 39'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_pc <= 39'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_pc <= frontend_io_out_0_bits_cf_pc;
            end else begin
              _T_6_1_cf_pc <= 39'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_pc <= frontend_io_out_0_bits_cf_pc;
          end else begin
            _T_6_1_cf_pc <= 39'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_pnpc <= 39'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_pnpc <= 39'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_pnpc <= frontend_io_out_0_bits_cf_pnpc;
            end else begin
              _T_6_1_cf_pnpc <= 39'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_pnpc <= frontend_io_out_0_bits_cf_pnpc;
          end else begin
            _T_6_1_cf_pnpc <= 39'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_exceptionVec_1 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_exceptionVec_1 <= 1'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            _T_6_1_cf_exceptionVec_1 <= _T_27_cf_exceptionVec_1;
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          _T_6_1_cf_exceptionVec_1 <= _T_27_cf_exceptionVec_1;
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_exceptionVec_2 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_exceptionVec_2 <= 1'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            _T_6_1_cf_exceptionVec_2 <= _T_27_cf_exceptionVec_2;
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          _T_6_1_cf_exceptionVec_2 <= _T_27_cf_exceptionVec_2;
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_exceptionVec_12 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_exceptionVec_12 <= 1'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            _T_6_1_cf_exceptionVec_12 <= _T_27_cf_exceptionVec_12;
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          _T_6_1_cf_exceptionVec_12 <= _T_27_cf_exceptionVec_12;
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_intrVec_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_intrVec_0 <= _T_6_T_29_cf_intrVec_0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_intrVec_0 <= frontend_io_out_0_bits_cf_intrVec_0;
            end else begin
              _T_6_1_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_intrVec_0 <= frontend_io_out_0_bits_cf_intrVec_0;
          end else begin
            _T_6_1_cf_intrVec_0 <= frontend_io_out_1_bits_cf_intrVec_0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_intrVec_1 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_intrVec_1 <= _T_6_T_29_cf_intrVec_1;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_intrVec_1 <= frontend_io_out_0_bits_cf_intrVec_1;
            end else begin
              _T_6_1_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_intrVec_1 <= frontend_io_out_0_bits_cf_intrVec_1;
          end else begin
            _T_6_1_cf_intrVec_1 <= frontend_io_out_1_bits_cf_intrVec_1;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_intrVec_2 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_intrVec_2 <= _T_6_T_29_cf_intrVec_2;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_intrVec_2 <= frontend_io_out_0_bits_cf_intrVec_2;
            end else begin
              _T_6_1_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_intrVec_2 <= frontend_io_out_0_bits_cf_intrVec_2;
          end else begin
            _T_6_1_cf_intrVec_2 <= frontend_io_out_1_bits_cf_intrVec_2;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_intrVec_3 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_intrVec_3 <= _T_6_T_29_cf_intrVec_3;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_intrVec_3 <= frontend_io_out_0_bits_cf_intrVec_3;
            end else begin
              _T_6_1_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_intrVec_3 <= frontend_io_out_0_bits_cf_intrVec_3;
          end else begin
            _T_6_1_cf_intrVec_3 <= frontend_io_out_1_bits_cf_intrVec_3;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_intrVec_4 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_intrVec_4 <= _T_6_T_29_cf_intrVec_4;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_intrVec_4 <= frontend_io_out_0_bits_cf_intrVec_4;
            end else begin
              _T_6_1_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_intrVec_4 <= frontend_io_out_0_bits_cf_intrVec_4;
          end else begin
            _T_6_1_cf_intrVec_4 <= frontend_io_out_1_bits_cf_intrVec_4;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_intrVec_5 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_intrVec_5 <= _T_6_T_29_cf_intrVec_5;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_intrVec_5 <= frontend_io_out_0_bits_cf_intrVec_5;
            end else begin
              _T_6_1_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_intrVec_5 <= frontend_io_out_0_bits_cf_intrVec_5;
          end else begin
            _T_6_1_cf_intrVec_5 <= frontend_io_out_1_bits_cf_intrVec_5;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_intrVec_6 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_intrVec_6 <= _T_6_T_29_cf_intrVec_6;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_intrVec_6 <= frontend_io_out_0_bits_cf_intrVec_6;
            end else begin
              _T_6_1_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_intrVec_6 <= frontend_io_out_0_bits_cf_intrVec_6;
          end else begin
            _T_6_1_cf_intrVec_6 <= frontend_io_out_1_bits_cf_intrVec_6;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_intrVec_7 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_intrVec_7 <= _T_6_T_29_cf_intrVec_7;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_intrVec_7 <= frontend_io_out_0_bits_cf_intrVec_7;
            end else begin
              _T_6_1_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_intrVec_7 <= frontend_io_out_0_bits_cf_intrVec_7;
          end else begin
            _T_6_1_cf_intrVec_7 <= frontend_io_out_1_bits_cf_intrVec_7;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_intrVec_8 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_intrVec_8 <= _T_6_T_29_cf_intrVec_8;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_intrVec_8 <= frontend_io_out_0_bits_cf_intrVec_8;
            end else begin
              _T_6_1_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_intrVec_8 <= frontend_io_out_0_bits_cf_intrVec_8;
          end else begin
            _T_6_1_cf_intrVec_8 <= frontend_io_out_1_bits_cf_intrVec_8;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_intrVec_9 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_intrVec_9 <= _T_6_T_29_cf_intrVec_9;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_intrVec_9 <= frontend_io_out_0_bits_cf_intrVec_9;
            end else begin
              _T_6_1_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_intrVec_9 <= frontend_io_out_0_bits_cf_intrVec_9;
          end else begin
            _T_6_1_cf_intrVec_9 <= frontend_io_out_1_bits_cf_intrVec_9;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_intrVec_10 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_intrVec_10 <= _T_6_T_29_cf_intrVec_10;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_intrVec_10 <= frontend_io_out_0_bits_cf_intrVec_10;
            end else begin
              _T_6_1_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_intrVec_10 <= frontend_io_out_0_bits_cf_intrVec_10;
          end else begin
            _T_6_1_cf_intrVec_10 <= frontend_io_out_1_bits_cf_intrVec_10;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_intrVec_11 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_intrVec_11 <= _T_6_T_29_cf_intrVec_11;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_intrVec_11 <= frontend_io_out_0_bits_cf_intrVec_11;
            end else begin
              _T_6_1_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_intrVec_11 <= frontend_io_out_0_bits_cf_intrVec_11;
          end else begin
            _T_6_1_cf_intrVec_11 <= frontend_io_out_1_bits_cf_intrVec_11;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_brIdx <= 4'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_brIdx <= 4'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_cf_brIdx <= frontend_io_out_0_bits_cf_brIdx;
            end else begin
              _T_6_1_cf_brIdx <= 4'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_cf_brIdx <= frontend_io_out_0_bits_cf_brIdx;
          end else begin
            _T_6_1_cf_brIdx <= 4'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_cf_crossPageIPFFix <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_cf_crossPageIPFFix <= 1'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            _T_6_1_cf_crossPageIPFFix <= _T_27_cf_crossPageIPFFix;
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          _T_6_1_cf_crossPageIPFFix <= _T_27_cf_crossPageIPFFix;
        end
      end
    end
    if (reset) begin
      _T_6_1_ctrl_src1Type <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        _T_6_1_ctrl_src1Type <= _GEN_485;
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_ctrl_src1Type <= frontend_io_out_0_bits_ctrl_src1Type;
          end else begin
            _T_6_1_ctrl_src1Type <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_ctrl_src2Type <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        _T_6_1_ctrl_src2Type <= _GEN_481;
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_ctrl_src2Type <= frontend_io_out_0_bits_ctrl_src2Type;
          end else begin
            _T_6_1_ctrl_src2Type <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_ctrl_fuType <= 3'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_ctrl_fuType <= 3'h3;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_ctrl_fuType <= frontend_io_out_0_bits_ctrl_fuType;
            end else begin
              _T_6_1_ctrl_fuType <= 3'h3;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_ctrl_fuType <= frontend_io_out_0_bits_ctrl_fuType;
          end else begin
            _T_6_1_ctrl_fuType <= 3'h3;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_ctrl_fuOpType <= 7'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_ctrl_fuOpType <= 7'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_ctrl_fuOpType <= frontend_io_out_0_bits_ctrl_fuOpType;
            end else begin
              _T_6_1_ctrl_fuOpType <= 7'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_ctrl_fuOpType <= frontend_io_out_0_bits_ctrl_fuOpType;
          end else begin
            _T_6_1_ctrl_fuOpType <= 7'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_ctrl_rfSrc1 <= 5'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_ctrl_rfSrc1 <= 5'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_ctrl_rfSrc1 <= frontend_io_out_0_bits_ctrl_rfSrc1;
            end else begin
              _T_6_1_ctrl_rfSrc1 <= 5'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_ctrl_rfSrc1 <= frontend_io_out_0_bits_ctrl_rfSrc1;
          end else begin
            _T_6_1_ctrl_rfSrc1 <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_ctrl_rfSrc2 <= 5'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_ctrl_rfSrc2 <= 5'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_ctrl_rfSrc2 <= frontend_io_out_0_bits_ctrl_rfSrc2;
            end else begin
              _T_6_1_ctrl_rfSrc2 <= 5'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_ctrl_rfSrc2 <= frontend_io_out_0_bits_ctrl_rfSrc2;
          end else begin
            _T_6_1_ctrl_rfSrc2 <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_ctrl_rfWen <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_ctrl_rfWen <= 1'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            _T_6_1_ctrl_rfWen <= _T_27_ctrl_rfWen;
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          _T_6_1_ctrl_rfWen <= _T_27_ctrl_rfWen;
        end
      end
    end
    if (reset) begin
      _T_6_1_ctrl_rfDest <= 5'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_ctrl_rfDest <= 5'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_ctrl_rfDest <= frontend_io_out_0_bits_ctrl_rfDest;
            end else begin
              _T_6_1_ctrl_rfDest <= 5'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_ctrl_rfDest <= frontend_io_out_0_bits_ctrl_rfDest;
          end else begin
            _T_6_1_ctrl_rfDest <= 5'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_1_data_imm <= 64'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h1 == _T_29) begin
          _T_6_1_data_imm <= 64'h0;
        end else if (_T_20) begin
          if (2'h1 == _T_25[1:0]) begin
            if (_T_18_0) begin
              _T_6_1_data_imm <= frontend_io_out_0_bits_data_imm;
            end else begin
              _T_6_1_data_imm <= 64'h0;
            end
          end
        end
      end else if (_T_20) begin
        if (2'h1 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_1_data_imm <= frontend_io_out_0_bits_data_imm;
          end else begin
            _T_6_1_data_imm <= 64'h0;
          end
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_instr <= 64'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_instr <= 64'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_instr <= _T_27_cf_instr;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_instr <= _T_27_cf_instr;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_pc <= 39'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_pc <= 39'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_pc <= _T_27_cf_pc;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_pc <= _T_27_cf_pc;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_pnpc <= 39'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_pnpc <= 39'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_pnpc <= _T_27_cf_pnpc;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_pnpc <= _T_27_cf_pnpc;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_exceptionVec_1 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_exceptionVec_1 <= 1'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_exceptionVec_1 <= _T_27_cf_exceptionVec_1;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_exceptionVec_1 <= _T_27_cf_exceptionVec_1;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_exceptionVec_2 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_exceptionVec_2 <= 1'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_exceptionVec_2 <= _T_27_cf_exceptionVec_2;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_exceptionVec_2 <= _T_27_cf_exceptionVec_2;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_exceptionVec_12 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_exceptionVec_12 <= 1'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_exceptionVec_12 <= _T_27_cf_exceptionVec_12;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_exceptionVec_12 <= _T_27_cf_exceptionVec_12;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_intrVec_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_intrVec_0 <= _T_6_T_29_cf_intrVec_0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_intrVec_0 <= _T_27_cf_intrVec_0;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_intrVec_0 <= _T_27_cf_intrVec_0;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_intrVec_1 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_intrVec_1 <= _T_6_T_29_cf_intrVec_1;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_intrVec_1 <= _T_27_cf_intrVec_1;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_intrVec_1 <= _T_27_cf_intrVec_1;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_intrVec_2 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_intrVec_2 <= _T_6_T_29_cf_intrVec_2;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_intrVec_2 <= _T_27_cf_intrVec_2;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_intrVec_2 <= _T_27_cf_intrVec_2;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_intrVec_3 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_intrVec_3 <= _T_6_T_29_cf_intrVec_3;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_intrVec_3 <= _T_27_cf_intrVec_3;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_intrVec_3 <= _T_27_cf_intrVec_3;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_intrVec_4 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_intrVec_4 <= _T_6_T_29_cf_intrVec_4;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_intrVec_4 <= _T_27_cf_intrVec_4;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_intrVec_4 <= _T_27_cf_intrVec_4;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_intrVec_5 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_intrVec_5 <= _T_6_T_29_cf_intrVec_5;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_intrVec_5 <= _T_27_cf_intrVec_5;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_intrVec_5 <= _T_27_cf_intrVec_5;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_intrVec_6 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_intrVec_6 <= _T_6_T_29_cf_intrVec_6;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_intrVec_6 <= _T_27_cf_intrVec_6;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_intrVec_6 <= _T_27_cf_intrVec_6;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_intrVec_7 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_intrVec_7 <= _T_6_T_29_cf_intrVec_7;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_intrVec_7 <= _T_27_cf_intrVec_7;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_intrVec_7 <= _T_27_cf_intrVec_7;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_intrVec_8 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_intrVec_8 <= _T_6_T_29_cf_intrVec_8;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_intrVec_8 <= _T_27_cf_intrVec_8;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_intrVec_8 <= _T_27_cf_intrVec_8;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_intrVec_9 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_intrVec_9 <= _T_6_T_29_cf_intrVec_9;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_intrVec_9 <= _T_27_cf_intrVec_9;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_intrVec_9 <= _T_27_cf_intrVec_9;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_intrVec_10 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_intrVec_10 <= _T_6_T_29_cf_intrVec_10;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_intrVec_10 <= _T_27_cf_intrVec_10;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_intrVec_10 <= _T_27_cf_intrVec_10;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_intrVec_11 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_intrVec_11 <= _T_6_T_29_cf_intrVec_11;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_intrVec_11 <= _T_27_cf_intrVec_11;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_intrVec_11 <= _T_27_cf_intrVec_11;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_brIdx <= 4'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_brIdx <= 4'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_brIdx <= _T_27_cf_brIdx;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_brIdx <= _T_27_cf_brIdx;
        end
      end
    end
    if (reset) begin
      _T_6_2_cf_crossPageIPFFix <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_cf_crossPageIPFFix <= 1'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_cf_crossPageIPFFix <= _T_27_cf_crossPageIPFFix;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_cf_crossPageIPFFix <= _T_27_cf_crossPageIPFFix;
        end
      end
    end
    if (reset) begin
      _T_6_2_ctrl_src1Type <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        _T_6_2_ctrl_src1Type <= _GEN_486;
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_2_ctrl_src1Type <= frontend_io_out_0_bits_ctrl_src1Type;
          end else begin
            _T_6_2_ctrl_src1Type <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_6_2_ctrl_src2Type <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        _T_6_2_ctrl_src2Type <= _GEN_482;
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_2_ctrl_src2Type <= frontend_io_out_0_bits_ctrl_src2Type;
          end else begin
            _T_6_2_ctrl_src2Type <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_6_2_ctrl_fuType <= 3'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_ctrl_fuType <= 3'h3;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_ctrl_fuType <= _T_27_ctrl_fuType;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_ctrl_fuType <= _T_27_ctrl_fuType;
        end
      end
    end
    if (reset) begin
      _T_6_2_ctrl_fuOpType <= 7'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_ctrl_fuOpType <= 7'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_ctrl_fuOpType <= _T_27_ctrl_fuOpType;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_ctrl_fuOpType <= _T_27_ctrl_fuOpType;
        end
      end
    end
    if (reset) begin
      _T_6_2_ctrl_rfSrc1 <= 5'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_ctrl_rfSrc1 <= 5'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_ctrl_rfSrc1 <= _T_27_ctrl_rfSrc1;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_ctrl_rfSrc1 <= _T_27_ctrl_rfSrc1;
        end
      end
    end
    if (reset) begin
      _T_6_2_ctrl_rfSrc2 <= 5'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_ctrl_rfSrc2 <= 5'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_ctrl_rfSrc2 <= _T_27_ctrl_rfSrc2;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_ctrl_rfSrc2 <= _T_27_ctrl_rfSrc2;
        end
      end
    end
    if (reset) begin
      _T_6_2_ctrl_rfWen <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_ctrl_rfWen <= 1'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_ctrl_rfWen <= _T_27_ctrl_rfWen;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_ctrl_rfWen <= _T_27_ctrl_rfWen;
        end
      end
    end
    if (reset) begin
      _T_6_2_ctrl_rfDest <= 5'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_ctrl_rfDest <= 5'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_ctrl_rfDest <= _T_27_ctrl_rfDest;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_ctrl_rfDest <= _T_27_ctrl_rfDest;
        end
      end
    end
    if (reset) begin
      _T_6_2_data_imm <= 64'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h2 == _T_29) begin
          _T_6_2_data_imm <= 64'h0;
        end else if (_T_20) begin
          if (2'h2 == _T_25[1:0]) begin
            _T_6_2_data_imm <= _T_27_data_imm;
          end
        end
      end else if (_T_20) begin
        if (2'h2 == _T_25[1:0]) begin
          _T_6_2_data_imm <= _T_27_data_imm;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_instr <= 64'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_instr <= 64'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_instr <= _T_27_cf_instr;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_instr <= _T_27_cf_instr;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_pc <= 39'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_pc <= 39'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_pc <= _T_27_cf_pc;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_pc <= _T_27_cf_pc;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_pnpc <= 39'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_pnpc <= 39'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_pnpc <= _T_27_cf_pnpc;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_pnpc <= _T_27_cf_pnpc;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_exceptionVec_1 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_exceptionVec_1 <= 1'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_exceptionVec_1 <= _T_27_cf_exceptionVec_1;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_exceptionVec_1 <= _T_27_cf_exceptionVec_1;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_exceptionVec_2 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_exceptionVec_2 <= 1'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_exceptionVec_2 <= _T_27_cf_exceptionVec_2;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_exceptionVec_2 <= _T_27_cf_exceptionVec_2;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_exceptionVec_12 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_exceptionVec_12 <= 1'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_exceptionVec_12 <= _T_27_cf_exceptionVec_12;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_exceptionVec_12 <= _T_27_cf_exceptionVec_12;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_intrVec_0 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_intrVec_0 <= _T_6_T_29_cf_intrVec_0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_intrVec_0 <= _T_27_cf_intrVec_0;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_intrVec_0 <= _T_27_cf_intrVec_0;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_intrVec_1 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_intrVec_1 <= _T_6_T_29_cf_intrVec_1;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_intrVec_1 <= _T_27_cf_intrVec_1;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_intrVec_1 <= _T_27_cf_intrVec_1;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_intrVec_2 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_intrVec_2 <= _T_6_T_29_cf_intrVec_2;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_intrVec_2 <= _T_27_cf_intrVec_2;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_intrVec_2 <= _T_27_cf_intrVec_2;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_intrVec_3 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_intrVec_3 <= _T_6_T_29_cf_intrVec_3;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_intrVec_3 <= _T_27_cf_intrVec_3;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_intrVec_3 <= _T_27_cf_intrVec_3;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_intrVec_4 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_intrVec_4 <= _T_6_T_29_cf_intrVec_4;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_intrVec_4 <= _T_27_cf_intrVec_4;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_intrVec_4 <= _T_27_cf_intrVec_4;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_intrVec_5 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_intrVec_5 <= _T_6_T_29_cf_intrVec_5;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_intrVec_5 <= _T_27_cf_intrVec_5;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_intrVec_5 <= _T_27_cf_intrVec_5;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_intrVec_6 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_intrVec_6 <= _T_6_T_29_cf_intrVec_6;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_intrVec_6 <= _T_27_cf_intrVec_6;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_intrVec_6 <= _T_27_cf_intrVec_6;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_intrVec_7 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_intrVec_7 <= _T_6_T_29_cf_intrVec_7;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_intrVec_7 <= _T_27_cf_intrVec_7;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_intrVec_7 <= _T_27_cf_intrVec_7;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_intrVec_8 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_intrVec_8 <= _T_6_T_29_cf_intrVec_8;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_intrVec_8 <= _T_27_cf_intrVec_8;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_intrVec_8 <= _T_27_cf_intrVec_8;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_intrVec_9 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_intrVec_9 <= _T_6_T_29_cf_intrVec_9;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_intrVec_9 <= _T_27_cf_intrVec_9;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_intrVec_9 <= _T_27_cf_intrVec_9;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_intrVec_10 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_intrVec_10 <= _T_6_T_29_cf_intrVec_10;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_intrVec_10 <= _T_27_cf_intrVec_10;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_intrVec_10 <= _T_27_cf_intrVec_10;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_intrVec_11 <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_intrVec_11 <= _T_6_T_29_cf_intrVec_11;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_intrVec_11 <= _T_27_cf_intrVec_11;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_intrVec_11 <= _T_27_cf_intrVec_11;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_brIdx <= 4'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_brIdx <= 4'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_brIdx <= _T_27_cf_brIdx;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_brIdx <= _T_27_cf_brIdx;
        end
      end
    end
    if (reset) begin
      _T_6_3_cf_crossPageIPFFix <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_cf_crossPageIPFFix <= 1'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_cf_crossPageIPFFix <= _T_27_cf_crossPageIPFFix;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_cf_crossPageIPFFix <= _T_27_cf_crossPageIPFFix;
        end
      end
    end
    if (reset) begin
      _T_6_3_ctrl_src1Type <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        _T_6_3_ctrl_src1Type <= _GEN_487;
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_3_ctrl_src1Type <= frontend_io_out_0_bits_ctrl_src1Type;
          end else begin
            _T_6_3_ctrl_src1Type <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_6_3_ctrl_src2Type <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        _T_6_3_ctrl_src2Type <= _GEN_483;
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          if (_T_18_0) begin
            _T_6_3_ctrl_src2Type <= frontend_io_out_0_bits_ctrl_src2Type;
          end else begin
            _T_6_3_ctrl_src2Type <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_6_3_ctrl_fuType <= 3'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_ctrl_fuType <= 3'h3;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_ctrl_fuType <= _T_27_ctrl_fuType;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_ctrl_fuType <= _T_27_ctrl_fuType;
        end
      end
    end
    if (reset) begin
      _T_6_3_ctrl_fuOpType <= 7'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_ctrl_fuOpType <= 7'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_ctrl_fuOpType <= _T_27_ctrl_fuOpType;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_ctrl_fuOpType <= _T_27_ctrl_fuOpType;
        end
      end
    end
    if (reset) begin
      _T_6_3_ctrl_rfSrc1 <= 5'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_ctrl_rfSrc1 <= 5'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_ctrl_rfSrc1 <= _T_27_ctrl_rfSrc1;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_ctrl_rfSrc1 <= _T_27_ctrl_rfSrc1;
        end
      end
    end
    if (reset) begin
      _T_6_3_ctrl_rfSrc2 <= 5'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_ctrl_rfSrc2 <= 5'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_ctrl_rfSrc2 <= _T_27_ctrl_rfSrc2;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_ctrl_rfSrc2 <= _T_27_ctrl_rfSrc2;
        end
      end
    end
    if (reset) begin
      _T_6_3_ctrl_rfWen <= 1'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_ctrl_rfWen <= 1'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_ctrl_rfWen <= _T_27_ctrl_rfWen;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_ctrl_rfWen <= _T_27_ctrl_rfWen;
        end
      end
    end
    if (reset) begin
      _T_6_3_ctrl_rfDest <= 5'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_ctrl_rfDest <= 5'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_ctrl_rfDest <= _T_27_ctrl_rfDest;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_ctrl_rfDest <= _T_27_ctrl_rfDest;
        end
      end
    end
    if (reset) begin
      _T_6_3_data_imm <= 64'h0;
    end else if (_T_22) begin
      if (_T_21) begin
        if (2'h3 == _T_29) begin
          _T_6_3_data_imm <= 64'h0;
        end else if (_T_20) begin
          if (2'h3 == _T_25[1:0]) begin
            _T_6_3_data_imm <= _T_27_data_imm;
          end
        end
      end else if (_T_20) begin
        if (2'h3 == _T_25[1:0]) begin
          _T_6_3_data_imm <= _T_27_data_imm;
        end
      end
    end
    if (reset) begin
      _T_7 <= 2'h0;
    end else if (frontend_io_flushVec[1]) begin
      _T_7 <= 2'h0;
    end else if (_T_22) begin
      _T_7 <= _T_31;
    end
    if (reset) begin
      _T_8 <= 2'h0;
    end else if (frontend_io_flushVec[1]) begin
      _T_8 <= 2'h0;
    end else if (_T_44) begin
      _T_8 <= _T_46;
    end
  end
endmodule
module CoherenceManager(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [3:0]  io_in_req_bits_cmd,
  input  [63:0] io_in_req_bits_wdata,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_mem_req_ready,
  output        io_out_mem_req_valid,
  output [31:0] io_out_mem_req_bits_addr,
  output [3:0]  io_out_mem_req_bits_cmd,
  output [63:0] io_out_mem_req_bits_wdata,
  output        io_out_mem_resp_ready,
  input         io_out_mem_resp_valid,
  input  [3:0]  io_out_mem_resp_bits_cmd,
  input  [63:0] io_out_mem_resp_bits_rdata,
  input         io_out_coh_req_ready,
  output        io_out_coh_req_valid,
  output [31:0] io_out_coh_req_bits_addr,
  output [63:0] io_out_coh_req_bits_wdata,
  output        io_out_coh_resp_ready,
  input         io_out_coh_resp_valid,
  input  [3:0]  io_out_coh_resp_bits_cmd,
  input  [63:0] io_out_coh_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [63:0] _RAND_3;
`endif // RANDOMIZE_REG_INIT
  reg [2:0] state; // @[Coherence.scala 45:22]
  wire  inflight = state != 3'h0; // @[Coherence.scala 46:24]
  wire  _T_1 = ~io_in_req_bits_cmd[0]; // @[SimpleBus.scala 73:18]
  wire  _T_3 = ~io_in_req_bits_cmd[3]; // @[SimpleBus.scala 73:29]
  wire  _T_4 = _T_1 & _T_3; // @[SimpleBus.scala 73:26]
  wire  _T_5 = ~_T_4; // @[Coherence.scala 49:29]
  wire  _T_6 = io_in_req_valid & _T_5; // @[Coherence.scala 49:26]
  wire  _T_9 = _T_6 & _T_1; // @[Coherence.scala 49:52]
  wire  _T_10 = ~_T_9; // @[Coherence.scala 49:10]
  wire  _T_12 = _T_10 | reset; // @[Coherence.scala 49:9]
  wire  _T_13 = ~_T_12; // @[Coherence.scala 49:9]
  wire  _T_14 = ~inflight; // @[Coherence.scala 52:42]
  wire  _T_20 = _T_14 & _T_4; // @[Coherence.scala 52:52]
  reg [31:0] reqLatch_addr; // @[Reg.scala 15:16]
  reg [3:0] reqLatch_cmd; // @[Reg.scala 15:16]
  reg [63:0] reqLatch_wdata; // @[Reg.scala 15:16]
  wire  _T_23 = io_in_req_valid & _T_14; // @[Coherence.scala 65:43]
  wire  _T_25 = io_out_mem_req_ready & _T_14; // @[Coherence.scala 66:43]
  wire  _T_34 = io_out_coh_req_ready & _T_14; // @[Coherence.scala 69:43]
  wire  _GEN_5 = _T_4 & _T_23; // @[Coherence.scala 67:39]
  wire  _GEN_6 = _T_4 & _T_34; // @[Coherence.scala 67:39]
  wire  _GEN_7 = io_in_req_bits_cmd[0] & _T_23; // @[Coherence.scala 64:61]
  wire  _T_35 = 3'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_36 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_43 = io_in_req_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_44 = 3'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_45 = io_out_coh_resp_ready & io_out_coh_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_46 = io_out_coh_resp_bits_cmd == 4'hc; // @[SimpleBus.scala 92:26]
  wire  _T_48 = 3'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_50 = io_in_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire  _T_51 = io_in_resp_valid & _T_50; // @[Coherence.scala 89:29]
  wire  _T_52 = 3'h3 == state; // @[Conditional.scala 37:30]
  wire  _T_53 = io_out_mem_req_ready & io_out_mem_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_54 = 3'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_55 = io_out_mem_resp_ready & io_out_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_56 = io_out_mem_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire  _T_57 = _T_55 & _T_56; // @[Coherence.scala 96:55]
  wire  _T_58 = 3'h5 == state; // @[Conditional.scala 37:30]
  wire [63:0] _GEN_20 = _T_52 ? reqLatch_wdata : io_in_req_bits_wdata; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_22 = _T_52 ? reqLatch_cmd : io_in_req_bits_cmd; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_24 = _T_52 ? reqLatch_addr : io_in_req_bits_addr; // @[Conditional.scala 39:67]
  wire  _GEN_25 = _T_52 | _GEN_7; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_27 = _T_48 ? io_out_coh_resp_bits_rdata : io_out_mem_resp_bits_rdata; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_28 = _T_48 ? io_out_coh_resp_bits_cmd : io_out_mem_resp_bits_cmd; // @[Conditional.scala 39:67]
  wire  _GEN_29 = _T_48 ? io_out_coh_resp_valid : io_out_mem_resp_valid; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_32 = _T_48 ? io_in_req_bits_wdata : _GEN_20; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_34 = _T_48 ? io_in_req_bits_cmd : _GEN_22; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_36 = _T_48 ? io_in_req_bits_addr : _GEN_24; // @[Conditional.scala 39:67]
  wire  _GEN_37 = _T_48 ? _GEN_7 : _GEN_25; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_39 = _T_44 ? io_out_mem_resp_bits_rdata : _GEN_27; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_40 = _T_44 ? io_out_mem_resp_bits_cmd : _GEN_28; // @[Conditional.scala 39:67]
  wire  _GEN_41 = _T_44 ? io_out_mem_resp_valid : _GEN_29; // @[Conditional.scala 39:67]
  wire [63:0] _GEN_43 = _T_44 ? io_in_req_bits_wdata : _GEN_32; // @[Conditional.scala 39:67]
  wire [3:0] _GEN_45 = _T_44 ? io_in_req_bits_cmd : _GEN_34; // @[Conditional.scala 39:67]
  wire [31:0] _GEN_47 = _T_44 ? io_in_req_bits_addr : _GEN_36; // @[Conditional.scala 39:67]
  wire  _GEN_48 = _T_44 ? _GEN_7 : _GEN_37; // @[Conditional.scala 39:67]
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _T_25 : _GEN_6; // @[Coherence.scala 62:17 Coherence.scala 66:19 Coherence.scala 69:19]
  assign io_in_resp_valid = _T_35 ? io_out_mem_resp_valid : _GEN_41; // @[Coherence.scala 72:14 Coherence.scala 88:16]
  assign io_in_resp_bits_cmd = _T_35 ? io_out_mem_resp_bits_cmd : _GEN_40; // @[Coherence.scala 72:14 Coherence.scala 88:16]
  assign io_in_resp_bits_rdata = _T_35 ? io_out_mem_resp_bits_rdata : _GEN_39; // @[Coherence.scala 72:14 Coherence.scala 88:16]
  assign io_out_mem_req_valid = _T_35 ? _GEN_7 : _GEN_48; // @[Coherence.scala 61:24 Coherence.scala 65:26 Coherence.scala 93:28]
  assign io_out_mem_req_bits_addr = _T_35 ? io_in_req_bits_addr : _GEN_47; // @[Coherence.scala 59:23 Coherence.scala 92:27]
  assign io_out_mem_req_bits_cmd = _T_35 ? io_in_req_bits_cmd : _GEN_45; // @[Coherence.scala 59:23 Coherence.scala 92:27]
  assign io_out_mem_req_bits_wdata = _T_35 ? io_in_req_bits_wdata : _GEN_43; // @[Coherence.scala 59:23 Coherence.scala 92:27]
  assign io_out_mem_resp_ready = 1'h1; // @[Coherence.scala 72:14]
  assign io_out_coh_req_valid = io_in_req_bits_cmd[0] ? 1'h0 : _GEN_5; // @[Coherence.scala 63:24 Coherence.scala 68:26]
  assign io_out_coh_req_bits_addr = io_in_req_bits_addr; // @[Coherence.scala 54:16]
  assign io_out_coh_req_bits_wdata = io_in_req_bits_wdata; // @[Coherence.scala 54:16]
  assign io_out_coh_resp_ready = 1'h1; // @[Coherence.scala 56:18 Coherence.scala 88:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  reqLatch_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  reqLatch_cmd = _RAND_2[3:0];
  _RAND_3 = {2{`RANDOM}};
  reqLatch_wdata = _RAND_3[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 3'h0;
    end else if (_T_35) begin
      if (_T_36) begin
        if (_T_4) begin
          state <= 3'h1;
        end else if (_T_43) begin
          state <= 3'h5;
        end
      end
    end else if (_T_44) begin
      if (_T_45) begin
        if (_T_46) begin
          state <= 3'h2;
        end else begin
          state <= 3'h3;
        end
      end
    end else if (_T_48) begin
      if (_T_51) begin
        state <= 3'h0;
      end
    end else if (_T_52) begin
      if (_T_53) begin
        state <= 3'h4;
      end
    end else if (_T_54) begin
      if (_T_57) begin
        state <= 3'h0;
      end
    end else if (_T_58) begin
      if (_T_55) begin
        state <= 3'h0;
      end
    end
    if (_T_20) begin
      reqLatch_addr <= io_in_req_bits_addr;
    end
    if (_T_20) begin
      reqLatch_cmd <= io_in_req_bits_cmd;
    end
    if (_T_20) begin
      reqLatch_wdata <= io_in_req_bits_wdata;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_13) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Coherence.scala:49 assert(!(thisReq.valid && !thisReq.bits.isRead() && !thisReq.bits.isWrite()))\n"); // @[Coherence.scala 49:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_13) begin
          $fatal; // @[Coherence.scala 49:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module AXI42SimpleBusConverter(
  input         clock,
  input         reset,
  output        io_in_awready,
  input         io_in_awvalid,
  input  [31:0] io_in_awaddr,
  input  [17:0] io_in_awid,
  input  [7:0]  io_in_awlen,
  input  [2:0]  io_in_awsize,
  output        io_in_wready,
  input         io_in_wvalid,
  input  [63:0] io_in_wdata,
  input  [7:0]  io_in_wstrb,
  input         io_in_wlast,
  input         io_in_bready,
  output        io_in_bvalid,
  output        io_in_arready,
  input         io_in_arvalid,
  input  [31:0] io_in_araddr,
  input  [17:0] io_in_arid,
  input  [7:0]  io_in_arlen,
  input  [2:0]  io_in_arsize,
  input         io_in_rready,
  output        io_in_rvalid,
  output [63:0] io_in_rdata,
  output        io_in_rlast,
  output [17:0] io_in_rid,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [2:0]  io_out_req_bits_size,
  output [3:0]  io_out_req_bits_cmd,
  output [7:0]  io_out_req_bits_wmask,
  output [63:0] io_out_req_bits_wdata,
  output        io_out_resp_ready,
  input         io_out_resp_valid,
  input  [3:0]  io_out_resp_bits_cmd,
  input  [63:0] io_out_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg [17:0] inflight_id_reg; // @[ToAXI4.scala 38:32]
  reg [1:0] inflight_type; // @[ToAXI4.scala 40:30]
  wire  _T = inflight_type == 2'h0; // @[ToAXI4.scala 50:19]
  wire  _T_1 = ~_T; // @[ToAXI4.scala 53:5]
  wire  _T_2 = ~_T_1; // @[ToAXI4.scala 64:9]
  wire  _T_3 = _T_2 & io_in_arvalid; // @[ToAXI4.scala 64:23]
  wire  _T_4 = io_in_arlen == 8'h0; // @[ToAXI4.scala 67:27]
  wire [1:0] _T_5 = _T_4 ? 2'h0 : 2'h2; // @[ToAXI4.scala 67:19]
  wire  _T_6 = io_out_req_ready & io_out_req_valid; // @[Decoupled.scala 40:37]
  wire [31:0] _GEN_2 = _T_3 ? io_in_araddr : 32'h0; // @[ToAXI4.scala 64:40]
  wire [3:0] _GEN_3 = _T_3 ? {{2'd0}, _T_5} : 4'h0; // @[ToAXI4.scala 64:40]
  wire [2:0] _GEN_4 = _T_3 ? io_in_arsize : 3'h0; // @[ToAXI4.scala 64:40]
  wire  _T_7 = inflight_type == 2'h1; // @[ToAXI4.scala 50:19]
  wire  _T_8 = _T_7 & io_out_resp_valid; // @[ToAXI4.scala 79:27]
  wire  _T_9 = io_out_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire  _T_10 = io_in_rready & io_in_rvalid; // @[Decoupled.scala 40:37]
  wire  _T_12 = _T_10 & _T_9; // @[ToAXI4.scala 88:22]
  reg [31:0] aw_reg_addr; // @[ToAXI4.scala 94:19]
  reg [7:0] aw_reg_len; // @[ToAXI4.scala 94:19]
  reg [2:0] aw_reg_size; // @[ToAXI4.scala 94:19]
  reg  bresp_en; // @[ToAXI4.scala 95:25]
  wire  _T_16 = _T_2 & io_in_awvalid; // @[ToAXI4.scala 97:23]
  wire  _T_17 = ~io_in_arvalid; // @[ToAXI4.scala 97:42]
  wire  _T_18 = _T_16 & _T_17; // @[ToAXI4.scala 97:39]
  wire  _T_19 = io_in_awready & io_in_awvalid; // @[Decoupled.scala 40:37]
  wire  _T_20 = inflight_type == 2'h2; // @[ToAXI4.scala 50:19]
  wire  _T_21 = io_in_wready & io_in_wvalid; // @[Decoupled.scala 40:37]
  wire  _T_22 = _T_20 & _T_21; // @[ToAXI4.scala 105:28]
  wire  _T_23 = aw_reg_len == 8'h0; // @[ToAXI4.scala 107:31]
  wire [2:0] _T_24 = io_in_wlast ? 3'h7 : 3'h3; // @[ToAXI4.scala 108:10]
  wire [2:0] _T_25 = _T_23 ? 3'h1 : _T_24; // @[ToAXI4.scala 107:19]
  wire  _GEN_31 = io_in_wlast | bresp_en; // @[ToAXI4.scala 115:19]
  wire  _T_26 = io_in_bready & io_in_bvalid; // @[Decoupled.scala 40:37]
  wire  _T_32 = _T_20 & io_in_wvalid; // @[ToAXI4.scala 127:75]
  wire  _T_38 = _T_7 & io_in_rready; // @[ToAXI4.scala 128:57]
  wire  _T_39 = _T_2 | _T_38; // @[ToAXI4.scala 128:35]
  wire  _T_41 = _T_20 & io_in_bready; // @[ToAXI4.scala 128:96]
  wire  _T_57 = io_in_arready & io_in_arvalid; // @[Decoupled.scala 40:37]
  wire  _T_62 = _T_6 & _T_2; // @[ToAXI4.scala 137:48]
  wire  _T_64 = _T_62 | reset; // @[ToAXI4.scala 137:32]
  wire  _T_65 = ~_T_64; // @[ToAXI4.scala 137:32]
  wire  _T_71 = _T_2 | reset; // @[ToAXI4.scala 138:32]
  wire  _T_72 = ~_T_71; // @[ToAXI4.scala 138:32]
  wire  _T_76 = _T_6 & _T_20; // @[ToAXI4.scala 139:48]
  wire  _T_78 = _T_76 | reset; // @[ToAXI4.scala 139:31]
  wire  _T_79 = ~_T_78; // @[ToAXI4.scala 139:31]
  wire  _T_81 = io_out_resp_ready & io_out_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_83 = _T_81 & _T_20; // @[ToAXI4.scala 140:48]
  wire  _T_85 = _T_83 | reset; // @[ToAXI4.scala 140:31]
  wire  _T_86 = ~_T_85; // @[ToAXI4.scala 140:31]
  wire  _T_90 = _T_81 & _T_7; // @[ToAXI4.scala 141:48]
  wire  _T_92 = _T_90 | reset; // @[ToAXI4.scala 141:31]
  wire  _T_93 = ~_T_92; // @[ToAXI4.scala 141:31]
  assign io_in_awready = _T_2 & _T_17; // @[ToAXI4.scala 132:16]
  assign io_in_wready = _T_20 & io_out_req_ready; // @[ToAXI4.scala 133:16]
  assign io_in_bvalid = bresp_en & io_out_resp_valid; // @[ToAXI4.scala 134:15]
  assign io_in_arready = _T_2 & io_out_req_ready; // @[ToAXI4.scala 129:16]
  assign io_in_rvalid = _T_7 & io_out_resp_valid; // @[ToAXI4.scala 80:17 ToAXI4.scala 130:15]
  assign io_in_rdata = _T_8 ? io_out_resp_bits_rdata : 64'h0; // @[ToAXI4.scala 60:5 ToAXI4.scala 81:12]
  assign io_in_rlast = _T_8 & _T_9; // @[ToAXI4.scala 60:5 ToAXI4.scala 85:12]
  assign io_in_rid = _T_8 ? inflight_id_reg : 18'h0; // @[ToAXI4.scala 60:5 ToAXI4.scala 82:10]
  assign io_out_req_valid = _T_3 | _T_32; // @[ToAXI4.scala 65:19 ToAXI4.scala 106:19 ToAXI4.scala 127:17]
  assign io_out_req_bits_addr = _T_22 ? aw_reg_addr : _GEN_2; // @[ToAXI4.scala 59:7 ToAXI4.scala 66:14 ToAXI4.scala 109:14]
  assign io_out_req_bits_size = _T_22 ? aw_reg_size : _GEN_4; // @[ToAXI4.scala 59:7 ToAXI4.scala 69:14 ToAXI4.scala 110:14]
  assign io_out_req_bits_cmd = _T_22 ? {{1'd0}, _T_25} : _GEN_3; // @[ToAXI4.scala 59:7 ToAXI4.scala 67:13 ToAXI4.scala 107:13]
  assign io_out_req_bits_wmask = _T_22 ? io_in_wstrb : 8'h0; // @[ToAXI4.scala 59:7 ToAXI4.scala 71:15 ToAXI4.scala 111:15]
  assign io_out_req_bits_wdata = _T_22 ? io_in_wdata : 64'h0; // @[ToAXI4.scala 59:7 ToAXI4.scala 72:15 ToAXI4.scala 112:15]
  assign io_out_resp_ready = _T_39 | _T_41; // @[ToAXI4.scala 128:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inflight_id_reg = _RAND_0[17:0];
  _RAND_1 = {1{`RANDOM}};
  inflight_type = _RAND_1[1:0];
  _RAND_2 = {1{`RANDOM}};
  aw_reg_addr = _RAND_2[31:0];
  _RAND_3 = {1{`RANDOM}};
  aw_reg_len = _RAND_3[7:0];
  _RAND_4 = {1{`RANDOM}};
  aw_reg_size = _RAND_4[2:0];
  _RAND_5 = {1{`RANDOM}};
  bresp_en = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      inflight_id_reg <= 18'h0;
    end else if (_T_26) begin
      inflight_id_reg <= 18'h0;
    end else if (_T_18) begin
      if (_T_19) begin
        inflight_id_reg <= io_in_awid;
      end else if (_T_8) begin
        if (_T_12) begin
          inflight_id_reg <= 18'h0;
        end else if (_T_3) begin
          if (_T_6) begin
            inflight_id_reg <= io_in_arid;
          end
        end
      end else if (_T_3) begin
        if (_T_6) begin
          inflight_id_reg <= io_in_arid;
        end
      end
    end else if (_T_8) begin
      if (_T_12) begin
        inflight_id_reg <= 18'h0;
      end else if (_T_3) begin
        if (_T_6) begin
          inflight_id_reg <= io_in_arid;
        end
      end
    end else if (_T_3) begin
      if (_T_6) begin
        inflight_id_reg <= io_in_arid;
      end
    end
    if (reset) begin
      inflight_type <= 2'h0;
    end else if (_T_26) begin
      inflight_type <= 2'h0;
    end else if (_T_18) begin
      if (_T_19) begin
        inflight_type <= 2'h2;
      end else if (_T_8) begin
        if (_T_12) begin
          inflight_type <= 2'h0;
        end else if (_T_3) begin
          if (_T_6) begin
            inflight_type <= 2'h1;
          end
        end
      end else if (_T_3) begin
        if (_T_6) begin
          inflight_type <= 2'h1;
        end
      end
    end else if (_T_8) begin
      if (_T_12) begin
        inflight_type <= 2'h0;
      end else if (_T_3) begin
        if (_T_6) begin
          inflight_type <= 2'h1;
        end
      end
    end else if (_T_3) begin
      if (_T_6) begin
        inflight_type <= 2'h1;
      end
    end
    if (_T_18) begin
      aw_reg_addr <= io_in_awaddr;
    end
    if (_T_18) begin
      aw_reg_len <= io_in_awlen;
    end
    if (_T_18) begin
      aw_reg_size <= io_in_awsize;
    end
    if (reset) begin
      bresp_en <= 1'h0;
    end else if (_T_26) begin
      bresp_en <= 1'h0;
    end else if (_T_22) begin
      bresp_en <= _GEN_31;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_57 & _T_65) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:137 when (axi.ar.fire()) { assert(mem.req.fire() && !isInflight()); }\n"); // @[ToAXI4.scala 137:32]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_57 & _T_65) begin
          $fatal; // @[ToAXI4.scala 137:32]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_19 & _T_72) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:138 when (axi.aw.fire()) { assert(!isInflight()); }\n"); // @[ToAXI4.scala 138:32]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_19 & _T_72) begin
          $fatal; // @[ToAXI4.scala 138:32]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_21 & _T_79) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:139 when (axi.w.fire()) { assert(mem.req .fire() && isState(axi_write)); }\n"); // @[ToAXI4.scala 139:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_21 & _T_79) begin
          $fatal; // @[ToAXI4.scala 139:31]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_26 & _T_86) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:140 when (axi.b.fire()) { assert(mem.resp.fire() && isState(axi_write)); }\n"); // @[ToAXI4.scala 140:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_26 & _T_86) begin
          $fatal; // @[ToAXI4.scala 140:31]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_10 & _T_93) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:141 when (axi.r.fire()) { assert(mem.resp.fire() && isState(axi_read)); }\n"); // @[ToAXI4.scala 141:31]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_10 & _T_93) begin
          $fatal; // @[ToAXI4.scala 141:31]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Prefetcher(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [2:0]  io_in_bits_size,
  input  [3:0]  io_in_bits_cmd,
  input  [7:0]  io_in_bits_wmask,
  input  [63:0] io_in_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_addr,
  output [2:0]  io_out_bits_size,
  output [3:0]  io_out_bits_cmd,
  output [7:0]  io_out_bits_wmask,
  output [63:0] io_out_bits_wdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [63:0] _RAND_5;
`endif // RANDOMIZE_REG_INIT
  reg  getNewReq; // @[Prefetcher.scala 37:26]
  reg [31:0] prefetchReq_addr; // @[Prefetcher.scala 38:28]
  reg [2:0] prefetchReq_size; // @[Prefetcher.scala 38:28]
  reg [7:0] prefetchReq_wmask; // @[Prefetcher.scala 38:28]
  reg [63:0] prefetchReq_wdata; // @[Prefetcher.scala 38:28]
  reg [63:0] lastReqAddr; // @[Prefetcher.scala 44:28]
  wire  _T_2 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_9 = {{32'd0}, io_in_bits_addr}; // @[Prefetcher.scala 50:30]
  wire [63:0] _T_4 = _GEN_9 & 64'hffffffffffffffc0; // @[Prefetcher.scala 50:30]
  wire [63:0] _T_5 = lastReqAddr & 64'hffffffffffffffc0; // @[Prefetcher.scala 50:59]
  wire  neqAddr = _T_4 != _T_5; // @[Prefetcher.scala 50:42]
  wire  _T_6 = ~getNewReq; // @[Prefetcher.scala 52:9]
  wire  _T_7 = ~io_in_valid; // @[Prefetcher.scala 55:20]
  wire  _T_8 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_9 = _T_7 | _T_8; // @[Prefetcher.scala 55:33]
  wire  _T_12 = _T_2 & io_in_bits_cmd[1]; // @[Prefetcher.scala 56:31]
  wire  _T_13 = _T_12 & neqAddr; // @[Prefetcher.scala 56:55]
  wire [31:0] _T_14 = prefetchReq_addr ^ 32'h30000000; // @[NutCore.scala 86:11]
  wire  _T_16 = _T_14[31:28] == 4'h0; // @[NutCore.scala 86:44]
  wire [31:0] _T_17 = prefetchReq_addr ^ 32'he0000000; // @[NutCore.scala 86:11]
  wire  _T_19 = _T_17[31:29] == 3'h0; // @[NutCore.scala 86:44]
  wire  _T_20 = _T_16 | _T_19; // @[NutCore.scala 87:15]
  wire  _T_21 = ~_T_20; // @[Prefetcher.scala 59:21]
  wire  _T_30 = _T_8 | _T_20; // @[Prefetcher.scala 61:34]
  wire  _T_31 = ~_T_30; // @[Prefetcher.scala 61:18]
  assign io_in_ready = _T_6 & _T_9; // @[Prefetcher.scala 55:17 Prefetcher.scala 60:17]
  assign io_out_valid = _T_6 ? io_in_valid : _T_21; // @[Prefetcher.scala 54:18 Prefetcher.scala 59:18]
  assign io_out_bits_addr = _T_6 ? io_in_bits_addr : prefetchReq_addr; // @[Prefetcher.scala 53:17 Prefetcher.scala 58:17]
  assign io_out_bits_size = _T_6 ? io_in_bits_size : prefetchReq_size; // @[Prefetcher.scala 53:17 Prefetcher.scala 58:17]
  assign io_out_bits_cmd = _T_6 ? io_in_bits_cmd : 4'h4; // @[Prefetcher.scala 53:17 Prefetcher.scala 58:17]
  assign io_out_bits_wmask = _T_6 ? io_in_bits_wmask : prefetchReq_wmask; // @[Prefetcher.scala 53:17 Prefetcher.scala 58:17]
  assign io_out_bits_wdata = _T_6 ? io_in_bits_wdata : prefetchReq_wdata; // @[Prefetcher.scala 53:17 Prefetcher.scala 58:17]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  getNewReq = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  prefetchReq_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  prefetchReq_size = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  prefetchReq_wmask = _RAND_3[7:0];
  _RAND_4 = {2{`RANDOM}};
  prefetchReq_wdata = _RAND_4[63:0];
  _RAND_5 = {2{`RANDOM}};
  lastReqAddr = _RAND_5[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      getNewReq <= 1'h0;
    end else if (_T_6) begin
      getNewReq <= _T_13;
    end else begin
      getNewReq <= _T_31;
    end
    prefetchReq_addr <= io_in_bits_addr + 32'h40;
    prefetchReq_size <= io_in_bits_size;
    prefetchReq_wmask <= io_in_bits_wmask;
    prefetchReq_wdata <= io_in_bits_wdata;
    if (reset) begin
      lastReqAddr <= 64'h0;
    end else if (_T_2) begin
      lastReqAddr <= {{32'd0}, io_in_bits_addr};
    end
  end
endmodule
module CacheStage1_2(
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_addr,
  input  [3:0]  io_in_bits_cmd,
  input  [7:0]  io_in_bits_wmask,
  input  [63:0] io_in_bits_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [3:0]  io_out_bits_req_cmd,
  output [7:0]  io_out_bits_req_wmask,
  output [63:0] io_out_bits_req_wdata,
  input         io_metaReadBus_req_ready,
  output        io_metaReadBus_req_valid,
  output [8:0]  io_metaReadBus_req_bits_setIdx,
  input  [16:0] io_metaReadBus_resp_data_0_tag,
  input         io_metaReadBus_resp_data_0_valid,
  input         io_metaReadBus_resp_data_0_dirty,
  input  [16:0] io_metaReadBus_resp_data_1_tag,
  input         io_metaReadBus_resp_data_1_valid,
  input         io_metaReadBus_resp_data_1_dirty,
  input  [16:0] io_metaReadBus_resp_data_2_tag,
  input         io_metaReadBus_resp_data_2_valid,
  input         io_metaReadBus_resp_data_2_dirty,
  input  [16:0] io_metaReadBus_resp_data_3_tag,
  input         io_metaReadBus_resp_data_3_valid,
  input         io_metaReadBus_resp_data_3_dirty,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [11:0] io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data
);
  wire  _T_29 = io_in_valid & io_metaReadBus_req_ready; // @[Cache.scala 133:31]
  wire  _T_31 = ~io_in_valid; // @[Cache.scala 134:19]
  wire  _T_32 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  wire  _T_33 = _T_31 | _T_32; // @[Cache.scala 134:32]
  wire  _T_34 = _T_33 & io_metaReadBus_req_ready; // @[Cache.scala 134:50]
  assign io_in_ready = _T_34 & io_dataReadBus_req_ready; // @[Cache.scala 134:15]
  assign io_out_valid = _T_29 & io_dataReadBus_req_ready; // @[Cache.scala 133:16]
  assign io_out_bits_req_addr = io_in_bits_addr; // @[Cache.scala 132:19]
  assign io_out_bits_req_cmd = io_in_bits_cmd; // @[Cache.scala 132:19]
  assign io_out_bits_req_wmask = io_in_bits_wmask; // @[Cache.scala 132:19]
  assign io_out_bits_req_wdata = io_in_bits_wdata; // @[Cache.scala 132:19]
  assign io_metaReadBus_req_valid = io_in_valid & io_out_ready; // @[SRAMTemplate.scala 53:20]
  assign io_metaReadBus_req_bits_setIdx = io_in_bits_addr[14:6]; // @[SRAMTemplate.scala 26:17]
  assign io_dataReadBus_req_valid = io_in_valid & io_out_ready; // @[SRAMTemplate.scala 53:20]
  assign io_dataReadBus_req_bits_setIdx = {io_in_bits_addr[14:6],io_in_bits_addr[5:3]}; // @[SRAMTemplate.scala 26:17]
endmodule
module CacheStage2_2(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [3:0]  io_in_bits_req_cmd,
  input  [7:0]  io_in_bits_req_wmask,
  input  [63:0] io_in_bits_req_wdata,
  input         io_out_ready,
  output        io_out_valid,
  output [31:0] io_out_bits_req_addr,
  output [3:0]  io_out_bits_req_cmd,
  output [7:0]  io_out_bits_req_wmask,
  output [63:0] io_out_bits_req_wdata,
  output [16:0] io_out_bits_metas_0_tag,
  output        io_out_bits_metas_0_valid,
  output        io_out_bits_metas_0_dirty,
  output [16:0] io_out_bits_metas_1_tag,
  output        io_out_bits_metas_1_valid,
  output        io_out_bits_metas_1_dirty,
  output [16:0] io_out_bits_metas_2_tag,
  output        io_out_bits_metas_2_valid,
  output        io_out_bits_metas_2_dirty,
  output [16:0] io_out_bits_metas_3_tag,
  output        io_out_bits_metas_3_valid,
  output        io_out_bits_metas_3_dirty,
  output [63:0] io_out_bits_datas_0_data,
  output [63:0] io_out_bits_datas_1_data,
  output [63:0] io_out_bits_datas_2_data,
  output [63:0] io_out_bits_datas_3_data,
  output        io_out_bits_hit,
  output [3:0]  io_out_bits_waymask,
  output        io_out_bits_mmio,
  output        io_out_bits_isForwardData,
  output [63:0] io_out_bits_forwardData_data_data,
  output [3:0]  io_out_bits_forwardData_waymask,
  input  [16:0] io_metaReadResp_0_tag,
  input         io_metaReadResp_0_valid,
  input         io_metaReadResp_0_dirty,
  input  [16:0] io_metaReadResp_1_tag,
  input         io_metaReadResp_1_valid,
  input         io_metaReadResp_1_dirty,
  input  [16:0] io_metaReadResp_2_tag,
  input         io_metaReadResp_2_valid,
  input         io_metaReadResp_2_dirty,
  input  [16:0] io_metaReadResp_3_tag,
  input         io_metaReadResp_3_valid,
  input         io_metaReadResp_3_dirty,
  input  [63:0] io_dataReadResp_0_data,
  input  [63:0] io_dataReadResp_1_data,
  input  [63:0] io_dataReadResp_2_data,
  input  [63:0] io_dataReadResp_3_data,
  input         io_metaWriteBus_req_valid,
  input  [8:0]  io_metaWriteBus_req_bits_setIdx,
  input  [16:0] io_metaWriteBus_req_bits_data_tag,
  input         io_metaWriteBus_req_bits_data_dirty,
  input  [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_dataWriteBus_req_valid,
  input  [11:0] io_dataWriteBus_req_bits_setIdx,
  input  [63:0] io_dataWriteBus_req_bits_data_data,
  input  [3:0]  io_dataWriteBus_req_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [31:0] _RAND_7;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 162:31]
  wire [8:0] addr_index = io_in_bits_req_addr[14:6]; // @[Cache.scala 162:31]
  wire [16:0] addr_tag = io_in_bits_req_addr[31:15]; // @[Cache.scala 162:31]
  wire  _T_5 = io_in_valid & io_metaWriteBus_req_valid; // @[Cache.scala 164:35]
  wire  _T_12 = io_metaWriteBus_req_bits_setIdx == addr_index; // @[Cache.scala 164:99]
  wire  isForwardMeta = _T_5 & _T_12; // @[Cache.scala 164:64]
  reg  isForwardMetaReg; // @[Cache.scala 165:33]
  wire  _GEN_0 = isForwardMeta | isForwardMetaReg; // @[Cache.scala 166:24]
  wire  _T_13 = io_in_ready & io_in_valid; // @[Decoupled.scala 40:37]
  wire  _T_14 = ~io_in_valid; // @[Cache.scala 167:25]
  wire  _T_15 = _T_13 | _T_14; // @[Cache.scala 167:22]
  reg [16:0] forwardMetaReg_data_tag; // @[Reg.scala 15:16]
  reg  forwardMetaReg_data_dirty; // @[Reg.scala 15:16]
  reg [3:0] forwardMetaReg_waymask; // @[Reg.scala 15:16]
  wire [3:0] _GEN_2 = isForwardMeta ? io_metaWriteBus_req_bits_waymask : forwardMetaReg_waymask; // @[Reg.scala 16:19]
  wire  _GEN_3 = isForwardMeta ? io_metaWriteBus_req_bits_data_dirty : forwardMetaReg_data_dirty; // @[Reg.scala 16:19]
  wire [16:0] _GEN_5 = isForwardMeta ? io_metaWriteBus_req_bits_data_tag : forwardMetaReg_data_tag; // @[Reg.scala 16:19]
  wire  pickForwardMeta = isForwardMetaReg | isForwardMeta; // @[Cache.scala 171:42]
  wire  forwardWaymask_0 = _GEN_2[0]; // @[Cache.scala 173:61]
  wire  forwardWaymask_1 = _GEN_2[1]; // @[Cache.scala 173:61]
  wire  forwardWaymask_2 = _GEN_2[2]; // @[Cache.scala 173:61]
  wire  forwardWaymask_3 = _GEN_2[3]; // @[Cache.scala 173:61]
  wire  _T_16 = pickForwardMeta & forwardWaymask_0; // @[Cache.scala 175:39]
  wire [16:0] metaWay_0_tag = _T_16 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 175:22]
  wire  metaWay_0_valid = _T_16 | io_metaReadResp_0_valid; // @[Cache.scala 175:22]
  wire  _T_18 = pickForwardMeta & forwardWaymask_1; // @[Cache.scala 175:39]
  wire [16:0] metaWay_1_tag = _T_18 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 175:22]
  wire  metaWay_1_valid = _T_18 | io_metaReadResp_1_valid; // @[Cache.scala 175:22]
  wire  _T_20 = pickForwardMeta & forwardWaymask_2; // @[Cache.scala 175:39]
  wire [16:0] metaWay_2_tag = _T_20 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 175:22]
  wire  metaWay_2_valid = _T_20 | io_metaReadResp_2_valid; // @[Cache.scala 175:22]
  wire  _T_22 = pickForwardMeta & forwardWaymask_3; // @[Cache.scala 175:39]
  wire [16:0] metaWay_3_tag = _T_22 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 175:22]
  wire  metaWay_3_valid = _T_22 | io_metaReadResp_3_valid; // @[Cache.scala 175:22]
  wire  _T_24 = metaWay_0_tag == addr_tag; // @[Cache.scala 178:59]
  wire  _T_25 = metaWay_0_valid & _T_24; // @[Cache.scala 178:49]
  wire  _T_26 = _T_25 & io_in_valid; // @[Cache.scala 178:73]
  wire  _T_27 = metaWay_1_tag == addr_tag; // @[Cache.scala 178:59]
  wire  _T_28 = metaWay_1_valid & _T_27; // @[Cache.scala 178:49]
  wire  _T_29 = _T_28 & io_in_valid; // @[Cache.scala 178:73]
  wire  _T_30 = metaWay_2_tag == addr_tag; // @[Cache.scala 178:59]
  wire  _T_31 = metaWay_2_valid & _T_30; // @[Cache.scala 178:49]
  wire  _T_32 = _T_31 & io_in_valid; // @[Cache.scala 178:73]
  wire  _T_33 = metaWay_3_tag == addr_tag; // @[Cache.scala 178:59]
  wire  _T_34 = metaWay_3_valid & _T_33; // @[Cache.scala 178:49]
  wire  _T_35 = _T_34 & io_in_valid; // @[Cache.scala 178:73]
  wire [3:0] hitVec = {_T_35,_T_32,_T_29,_T_26}; // @[Cache.scala 178:90]
  reg [63:0] _T_39; // @[LFSR64.scala 25:23]
  wire  _T_42 = _T_39[0] ^ _T_39[1]; // @[LFSR64.scala 26:23]
  wire  _T_44 = _T_42 ^ _T_39[3]; // @[LFSR64.scala 26:33]
  wire  _T_46 = _T_44 ^ _T_39[4]; // @[LFSR64.scala 26:43]
  wire  _T_47 = _T_39 == 64'h0; // @[LFSR64.scala 28:24]
  wire [63:0] _T_49 = {_T_46,_T_39[63:1]}; // @[Cat.scala 29:58]
  wire [3:0] victimWaymask = 4'h1 << _T_39[1:0]; // @[Cache.scala 179:42]
  wire  _T_52 = ~metaWay_0_valid; // @[Cache.scala 181:45]
  wire  _T_53 = ~metaWay_1_valid; // @[Cache.scala 181:45]
  wire  _T_54 = ~metaWay_2_valid; // @[Cache.scala 181:45]
  wire  _T_55 = ~metaWay_3_valid; // @[Cache.scala 181:45]
  wire [3:0] invalidVec = {_T_55,_T_54,_T_53,_T_52}; // @[Cache.scala 181:56]
  wire  hasInvalidWay = |invalidVec; // @[Cache.scala 182:34]
  wire  _T_59 = invalidVec >= 4'h8; // @[Cache.scala 183:45]
  wire  _T_60 = invalidVec >= 4'h4; // @[Cache.scala 184:20]
  wire  _T_61 = invalidVec >= 4'h2; // @[Cache.scala 185:20]
  wire [1:0] _T_62 = _T_61 ? 2'h2 : 2'h1; // @[Cache.scala 185:8]
  wire [2:0] _T_63 = _T_60 ? 3'h4 : {{1'd0}, _T_62}; // @[Cache.scala 184:8]
  wire [3:0] refillInvalidWaymask = _T_59 ? 4'h8 : {{1'd0}, _T_63}; // @[Cache.scala 183:33]
  wire [3:0] _T_64 = hasInvalidWay ? refillInvalidWaymask : victimWaymask; // @[Cache.scala 188:49]
  wire [3:0] waymask = io_out_bits_hit ? hitVec : _T_64; // @[Cache.scala 188:20]
  wire [1:0] _T_69 = waymask[0] + waymask[1]; // @[Bitwise.scala 47:55]
  wire [1:0] _T_71 = waymask[2] + waymask[3]; // @[Bitwise.scala 47:55]
  wire [2:0] _T_73 = _T_69 + _T_71; // @[Bitwise.scala 47:55]
  wire  _T_75 = _T_73 > 3'h1; // @[Cache.scala 189:26]
  wire  _T_197 = io_in_valid & _T_75; // @[Cache.scala 196:24]
  wire  _T_198 = ~_T_197; // @[Cache.scala 196:10]
  wire  _T_200 = _T_198 | reset; // @[Cache.scala 196:9]
  wire  _T_201 = ~_T_200; // @[Cache.scala 196:9]
  wire  _T_202 = |hitVec; // @[Cache.scala 199:44]
  wire [31:0] _T_204 = io_in_bits_req_addr ^ 32'h30000000; // @[NutCore.scala 86:11]
  wire  _T_206 = _T_204[31:28] == 4'h0; // @[NutCore.scala 86:44]
  wire [31:0] _T_207 = io_in_bits_req_addr ^ 32'he0000000; // @[NutCore.scala 86:11]
  wire  _T_209 = _T_207[31:29] == 3'h0; // @[NutCore.scala 86:44]
  wire [11:0] _T_223 = {addr_index,addr_wordIndex}; // @[Cat.scala 29:58]
  wire  _T_224 = io_dataWriteBus_req_bits_setIdx == _T_223; // @[Cache.scala 205:30]
  wire  _T_225 = io_dataWriteBus_req_valid & _T_224; // @[Cache.scala 205:13]
  wire  isForwardData = io_in_valid & _T_225; // @[Cache.scala 204:35]
  reg  isForwardDataReg; // @[Cache.scala 207:33]
  wire  _GEN_8 = isForwardData | isForwardDataReg; // @[Cache.scala 208:24]
  reg [63:0] forwardDataReg_data_data; // @[Reg.scala 15:16]
  reg [3:0] forwardDataReg_waymask; // @[Reg.scala 15:16]
  wire  _T_232 = io_out_ready & io_out_valid; // @[Decoupled.scala 40:37]
  assign io_in_ready = _T_14 | _T_232; // @[Cache.scala 216:15]
  assign io_out_valid = io_in_valid; // @[Cache.scala 215:16]
  assign io_out_bits_req_addr = io_in_bits_req_addr; // @[Cache.scala 214:19]
  assign io_out_bits_req_cmd = io_in_bits_req_cmd; // @[Cache.scala 214:19]
  assign io_out_bits_req_wmask = io_in_bits_req_wmask; // @[Cache.scala 214:19]
  assign io_out_bits_req_wdata = io_in_bits_req_wdata; // @[Cache.scala 214:19]
  assign io_out_bits_metas_0_tag = _T_16 ? _GEN_5 : io_metaReadResp_0_tag; // @[Cache.scala 198:21]
  assign io_out_bits_metas_0_valid = _T_16 | io_metaReadResp_0_valid; // @[Cache.scala 198:21]
  assign io_out_bits_metas_0_dirty = _T_16 ? _GEN_3 : io_metaReadResp_0_dirty; // @[Cache.scala 198:21]
  assign io_out_bits_metas_1_tag = _T_18 ? _GEN_5 : io_metaReadResp_1_tag; // @[Cache.scala 198:21]
  assign io_out_bits_metas_1_valid = _T_18 | io_metaReadResp_1_valid; // @[Cache.scala 198:21]
  assign io_out_bits_metas_1_dirty = _T_18 ? _GEN_3 : io_metaReadResp_1_dirty; // @[Cache.scala 198:21]
  assign io_out_bits_metas_2_tag = _T_20 ? _GEN_5 : io_metaReadResp_2_tag; // @[Cache.scala 198:21]
  assign io_out_bits_metas_2_valid = _T_20 | io_metaReadResp_2_valid; // @[Cache.scala 198:21]
  assign io_out_bits_metas_2_dirty = _T_20 ? _GEN_3 : io_metaReadResp_2_dirty; // @[Cache.scala 198:21]
  assign io_out_bits_metas_3_tag = _T_22 ? _GEN_5 : io_metaReadResp_3_tag; // @[Cache.scala 198:21]
  assign io_out_bits_metas_3_valid = _T_22 | io_metaReadResp_3_valid; // @[Cache.scala 198:21]
  assign io_out_bits_metas_3_dirty = _T_22 ? _GEN_3 : io_metaReadResp_3_dirty; // @[Cache.scala 198:21]
  assign io_out_bits_datas_0_data = io_dataReadResp_0_data; // @[Cache.scala 201:21]
  assign io_out_bits_datas_1_data = io_dataReadResp_1_data; // @[Cache.scala 201:21]
  assign io_out_bits_datas_2_data = io_dataReadResp_2_data; // @[Cache.scala 201:21]
  assign io_out_bits_datas_3_data = io_dataReadResp_3_data; // @[Cache.scala 201:21]
  assign io_out_bits_hit = io_in_valid & _T_202; // @[Cache.scala 199:19]
  assign io_out_bits_waymask = io_out_bits_hit ? hitVec : _T_64; // @[Cache.scala 200:23]
  assign io_out_bits_mmio = _T_206 | _T_209; // @[Cache.scala 202:20]
  assign io_out_bits_isForwardData = isForwardDataReg | isForwardData; // @[Cache.scala 211:29]
  assign io_out_bits_forwardData_data_data = isForwardData ? io_dataWriteBus_req_bits_data_data : forwardDataReg_data_data; // @[Cache.scala 212:27]
  assign io_out_bits_forwardData_waymask = isForwardData ? io_dataWriteBus_req_bits_waymask : forwardDataReg_waymask; // @[Cache.scala 212:27]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  isForwardMetaReg = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  forwardMetaReg_data_tag = _RAND_1[16:0];
  _RAND_2 = {1{`RANDOM}};
  forwardMetaReg_data_dirty = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  forwardMetaReg_waymask = _RAND_3[3:0];
  _RAND_4 = {2{`RANDOM}};
  _T_39 = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  isForwardDataReg = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  forwardDataReg_data_data = _RAND_6[63:0];
  _RAND_7 = {1{`RANDOM}};
  forwardDataReg_waymask = _RAND_7[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      isForwardMetaReg <= 1'h0;
    end else if (_T_15) begin
      isForwardMetaReg <= 1'h0;
    end else begin
      isForwardMetaReg <= _GEN_0;
    end
    if (isForwardMeta) begin
      forwardMetaReg_data_tag <= io_metaWriteBus_req_bits_data_tag;
    end
    if (isForwardMeta) begin
      forwardMetaReg_data_dirty <= io_metaWriteBus_req_bits_data_dirty;
    end
    if (isForwardMeta) begin
      forwardMetaReg_waymask <= io_metaWriteBus_req_bits_waymask;
    end
    if (reset) begin
      _T_39 <= 64'h1234567887654321;
    end else if (_T_47) begin
      _T_39 <= 64'h1;
    end else begin
      _T_39 <= _T_49;
    end
    if (reset) begin
      isForwardDataReg <= 1'h0;
    end else if (_T_15) begin
      isForwardDataReg <= 1'h0;
    end else begin
      isForwardDataReg <= _GEN_8;
    end
    if (isForwardData) begin
      forwardDataReg_data_data <= io_dataWriteBus_req_bits_data_data;
    end
    if (isForwardData) begin
      forwardDataReg_waymask <= io_dataWriteBus_req_bits_waymask;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_201) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Cache.scala:196 assert(!(io.in.valid && PopCount(waymask) > 1.U))\n"); // @[Cache.scala 196:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_201) begin
          $fatal; // @[Cache.scala 196:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Arbiter_10(
  input         io_in_0_valid,
  input  [8:0]  io_in_0_bits_setIdx,
  input  [16:0] io_in_0_bits_data_tag,
  input  [3:0]  io_in_0_bits_waymask,
  input         io_in_1_valid,
  input  [8:0]  io_in_1_bits_setIdx,
  input  [16:0] io_in_1_bits_data_tag,
  input         io_in_1_bits_data_dirty,
  input  [3:0]  io_in_1_bits_waymask,
  output        io_out_valid,
  output [8:0]  io_out_bits_setIdx,
  output [16:0] io_out_bits_data_tag,
  output        io_out_bits_data_dirty,
  output [3:0]  io_out_bits_waymask
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  _T_2 = ~grant_1; // @[Arbiter.scala 135:19]
  assign io_out_valid = _T_2 | io_in_1_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_data_tag = io_in_0_valid ? io_in_0_bits_data_tag : io_in_1_bits_data_tag; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_data_dirty = io_in_0_valid | io_in_1_bits_data_dirty; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_waymask = io_in_0_valid ? io_in_0_bits_waymask : io_in_1_bits_waymask; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
endmodule
module Arbiter_11(
  input         io_in_0_valid,
  input  [11:0] io_in_0_bits_setIdx,
  input  [63:0] io_in_0_bits_data_data,
  input  [3:0]  io_in_0_bits_waymask,
  input         io_in_1_valid,
  input  [11:0] io_in_1_bits_setIdx,
  input  [63:0] io_in_1_bits_data_data,
  input  [3:0]  io_in_1_bits_waymask,
  output        io_out_valid,
  output [11:0] io_out_bits_setIdx,
  output [63:0] io_out_bits_data_data,
  output [3:0]  io_out_bits_waymask
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  _T_2 = ~grant_1; // @[Arbiter.scala 135:19]
  assign io_out_valid = _T_2 | io_in_1_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_data_data = io_in_0_valid ? io_in_0_bits_data_data : io_in_1_bits_data_data; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
  assign io_out_bits_waymask = io_in_0_valid ? io_in_0_bits_waymask : io_in_1_bits_waymask; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
endmodule
module CacheStage3_2(
  input         clock,
  input         reset,
  output        io_in_ready,
  input         io_in_valid,
  input  [31:0] io_in_bits_req_addr,
  input  [3:0]  io_in_bits_req_cmd,
  input  [7:0]  io_in_bits_req_wmask,
  input  [63:0] io_in_bits_req_wdata,
  input  [16:0] io_in_bits_metas_0_tag,
  input         io_in_bits_metas_0_valid,
  input         io_in_bits_metas_0_dirty,
  input  [16:0] io_in_bits_metas_1_tag,
  input         io_in_bits_metas_1_valid,
  input         io_in_bits_metas_1_dirty,
  input  [16:0] io_in_bits_metas_2_tag,
  input         io_in_bits_metas_2_valid,
  input         io_in_bits_metas_2_dirty,
  input  [16:0] io_in_bits_metas_3_tag,
  input         io_in_bits_metas_3_valid,
  input         io_in_bits_metas_3_dirty,
  input  [63:0] io_in_bits_datas_0_data,
  input  [63:0] io_in_bits_datas_1_data,
  input  [63:0] io_in_bits_datas_2_data,
  input  [63:0] io_in_bits_datas_3_data,
  input         io_in_bits_hit,
  input  [3:0]  io_in_bits_waymask,
  input         io_in_bits_mmio,
  input         io_in_bits_isForwardData,
  input  [63:0] io_in_bits_forwardData_data_data,
  input  [3:0]  io_in_bits_forwardData_waymask,
  output        io_out_valid,
  output [3:0]  io_out_bits_cmd,
  output [63:0] io_out_bits_rdata,
  output        io_isFinish,
  input         io_dataReadBus_req_ready,
  output        io_dataReadBus_req_valid,
  output [11:0] io_dataReadBus_req_bits_setIdx,
  input  [63:0] io_dataReadBus_resp_data_0_data,
  input  [63:0] io_dataReadBus_resp_data_1_data,
  input  [63:0] io_dataReadBus_resp_data_2_data,
  input  [63:0] io_dataReadBus_resp_data_3_data,
  output        io_dataWriteBus_req_valid,
  output [11:0] io_dataWriteBus_req_bits_setIdx,
  output [63:0] io_dataWriteBus_req_bits_data_data,
  output [3:0]  io_dataWriteBus_req_bits_waymask,
  output        io_metaWriteBus_req_valid,
  output [8:0]  io_metaWriteBus_req_bits_setIdx,
  output [16:0] io_metaWriteBus_req_bits_data_tag,
  output        io_metaWriteBus_req_bits_data_dirty,
  output [3:0]  io_metaWriteBus_req_bits_waymask,
  input         io_mem_req_ready,
  output        io_mem_req_valid,
  output [31:0] io_mem_req_bits_addr,
  output [3:0]  io_mem_req_bits_cmd,
  output [63:0] io_mem_req_bits_wdata,
  output        io_mem_resp_ready,
  input         io_mem_resp_valid,
  input  [3:0]  io_mem_resp_bits_cmd,
  input  [63:0] io_mem_resp_bits_rdata,
  output        io_cohResp_valid,
  output        io_dataReadRespToL1
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [63:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
`endif // RANDOMIZE_REG_INIT
  wire  metaWriteArb_io_in_0_valid; // @[Cache.scala 241:28]
  wire [8:0] metaWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 241:28]
  wire [16:0] metaWriteArb_io_in_0_bits_data_tag; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_in_0_bits_waymask; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_in_1_valid; // @[Cache.scala 241:28]
  wire [8:0] metaWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 241:28]
  wire [16:0] metaWriteArb_io_in_1_bits_data_tag; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_in_1_bits_data_dirty; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_in_1_bits_waymask; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_out_valid; // @[Cache.scala 241:28]
  wire [8:0] metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 241:28]
  wire [16:0] metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 241:28]
  wire  metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 241:28]
  wire [3:0] metaWriteArb_io_out_bits_waymask; // @[Cache.scala 241:28]
  wire  dataWriteArb_io_in_0_valid; // @[Cache.scala 242:28]
  wire [11:0] dataWriteArb_io_in_0_bits_setIdx; // @[Cache.scala 242:28]
  wire [63:0] dataWriteArb_io_in_0_bits_data_data; // @[Cache.scala 242:28]
  wire [3:0] dataWriteArb_io_in_0_bits_waymask; // @[Cache.scala 242:28]
  wire  dataWriteArb_io_in_1_valid; // @[Cache.scala 242:28]
  wire [11:0] dataWriteArb_io_in_1_bits_setIdx; // @[Cache.scala 242:28]
  wire [63:0] dataWriteArb_io_in_1_bits_data_data; // @[Cache.scala 242:28]
  wire [3:0] dataWriteArb_io_in_1_bits_waymask; // @[Cache.scala 242:28]
  wire  dataWriteArb_io_out_valid; // @[Cache.scala 242:28]
  wire [11:0] dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 242:28]
  wire [63:0] dataWriteArb_io_out_bits_data_data; // @[Cache.scala 242:28]
  wire [3:0] dataWriteArb_io_out_bits_waymask; // @[Cache.scala 242:28]
  wire [2:0] addr_wordIndex = io_in_bits_req_addr[5:3]; // @[Cache.scala 245:31]
  wire [8:0] addr_index = io_in_bits_req_addr[14:6]; // @[Cache.scala 245:31]
  wire  mmio = io_in_valid & io_in_bits_mmio; // @[Cache.scala 246:26]
  wire  hit = io_in_valid & io_in_bits_hit; // @[Cache.scala 247:25]
  wire  _T_5 = ~io_in_bits_hit; // @[Cache.scala 248:29]
  wire  miss = io_in_valid & _T_5; // @[Cache.scala 248:26]
  wire  _T_7 = io_in_bits_req_cmd == 4'h8; // @[SimpleBus.scala 79:23]
  wire  probe = io_in_valid & _T_7; // @[Cache.scala 249:39]
  wire  _T_8 = io_in_bits_req_cmd == 4'h2; // @[SimpleBus.scala 76:27]
  wire  hitReadBurst = hit & _T_8; // @[Cache.scala 250:26]
  wire [18:0] _T_14 = {io_in_bits_metas_0_tag,io_in_bits_metas_0_valid,io_in_bits_metas_0_dirty}; // @[Mux.scala 27:72]
  wire [18:0] _T_15 = io_in_bits_waymask[0] ? _T_14 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_17 = {io_in_bits_metas_1_tag,io_in_bits_metas_1_valid,io_in_bits_metas_1_dirty}; // @[Mux.scala 27:72]
  wire [18:0] _T_18 = io_in_bits_waymask[1] ? _T_17 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_20 = {io_in_bits_metas_2_tag,io_in_bits_metas_2_valid,io_in_bits_metas_2_dirty}; // @[Mux.scala 27:72]
  wire [18:0] _T_21 = io_in_bits_waymask[2] ? _T_20 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_23 = {io_in_bits_metas_3_tag,io_in_bits_metas_3_valid,io_in_bits_metas_3_dirty}; // @[Mux.scala 27:72]
  wire [18:0] _T_24 = io_in_bits_waymask[3] ? _T_23 : 19'h0; // @[Mux.scala 27:72]
  wire [18:0] _T_25 = _T_15 | _T_18; // @[Mux.scala 27:72]
  wire [18:0] _T_26 = _T_25 | _T_21; // @[Mux.scala 27:72]
  wire [18:0] _T_27 = _T_26 | _T_24; // @[Mux.scala 27:72]
  wire  meta_dirty = _T_27[0]; // @[Mux.scala 27:72]
  wire [16:0] meta_tag = _T_27[18:2]; // @[Mux.scala 27:72]
  wire  _T_32 = mmio & hit; // @[Cache.scala 252:17]
  wire  _T_33 = ~_T_32; // @[Cache.scala 252:10]
  wire  _T_35 = _T_33 | reset; // @[Cache.scala 252:9]
  wire  _T_36 = ~_T_35; // @[Cache.scala 252:9]
  wire  _T_37 = io_in_bits_waymask == io_in_bits_forwardData_waymask; // @[Cache.scala 260:71]
  wire  useForwardData = io_in_bits_isForwardData & _T_37; // @[Cache.scala 260:49]
  wire [63:0] _T_42 = io_in_bits_waymask[0] ? io_in_bits_datas_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_43 = io_in_bits_waymask[1] ? io_in_bits_datas_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_44 = io_in_bits_waymask[2] ? io_in_bits_datas_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_45 = io_in_bits_waymask[3] ? io_in_bits_datas_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_46 = _T_42 | _T_43; // @[Mux.scala 27:72]
  wire [63:0] _T_47 = _T_46 | _T_44; // @[Mux.scala 27:72]
  wire [63:0] _T_48 = _T_47 | _T_45; // @[Mux.scala 27:72]
  wire [63:0] dataRead = useForwardData ? io_in_bits_forwardData_data_data : _T_48; // @[Cache.scala 262:21]
  wire [7:0] _T_64 = io_in_bits_req_wmask[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_66 = io_in_bits_req_wmask[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_68 = io_in_bits_req_wmask[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_70 = io_in_bits_req_wmask[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_72 = io_in_bits_req_wmask[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_74 = io_in_bits_req_wmask[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_76 = io_in_bits_req_wmask[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_78 = io_in_bits_req_wmask[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_85 = {_T_78,_T_76,_T_74,_T_72,_T_70,_T_68,_T_66,_T_64}; // @[Cat.scala 29:58]
  wire [63:0] wordMask = io_in_bits_req_cmd[0] ? _T_85 : 64'h0; // @[Cache.scala 263:21]
  reg [2:0] value; // @[Counter.scala 29:33]
  wire  _T_87 = io_in_bits_req_cmd == 4'h3; // @[Cache.scala 266:34]
  wire  _T_88 = io_in_bits_req_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_89 = _T_87 | _T_88; // @[Cache.scala 266:62]
  wire  _T_90 = io_out_valid & _T_89; // @[Cache.scala 266:22]
  wire [2:0] _T_93 = value + 3'h1; // @[Counter.scala 39:22]
  wire [2:0] _GEN_0 = _T_90 ? _T_93 : value; // @[Cache.scala 266:85]
  wire  hitWrite = hit & io_in_bits_req_cmd[0]; // @[Cache.scala 270:22]
  wire [63:0] _T_96 = io_in_bits_req_wdata & wordMask; // @[BitUtils.scala 32:13]
  wire [63:0] _T_97 = ~wordMask; // @[BitUtils.scala 32:38]
  wire [63:0] _T_98 = dataRead & _T_97; // @[BitUtils.scala 32:36]
  wire [2:0] _T_103 = _T_89 ? value : addr_wordIndex; // @[Cache.scala 273:51]
  wire  _T_105 = ~meta_dirty; // @[Cache.scala 276:25]
  wire  metaHitWriteBus_req_valid = hitWrite & _T_105; // @[Cache.scala 276:22]
  reg [3:0] state; // @[Cache.scala 281:22]
  reg [2:0] value_1; // @[Counter.scala 29:33]
  reg [2:0] value_2; // @[Counter.scala 29:33]
  reg [1:0] state2; // @[Cache.scala 291:23]
  wire  _T_118 = state == 4'h3; // @[Cache.scala 293:39]
  wire  _T_119 = state == 4'h8; // @[Cache.scala 293:66]
  wire  _T_120 = _T_118 | _T_119; // @[Cache.scala 293:57]
  wire  _T_121 = state2 == 2'h0; // @[Cache.scala 293:92]
  wire [2:0] _T_124 = _T_119 ? value_1 : value_2; // @[Cache.scala 294:33]
  wire  _T_126 = state2 == 2'h1; // @[Cache.scala 295:60]
  reg [63:0] dataWay_0_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_1_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_2_data; // @[Reg.scala 15:16]
  reg [63:0] dataWay_3_data; // @[Reg.scala 15:16]
  wire [63:0] _T_131 = io_in_bits_waymask[0] ? dataWay_0_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_132 = io_in_bits_waymask[1] ? dataWay_1_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_133 = io_in_bits_waymask[2] ? dataWay_2_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_134 = io_in_bits_waymask[3] ? dataWay_3_data : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_135 = _T_131 | _T_132; // @[Mux.scala 27:72]
  wire [63:0] _T_136 = _T_135 | _T_133; // @[Mux.scala 27:72]
  wire [63:0] _T_137 = _T_136 | _T_134; // @[Mux.scala 27:72]
  wire  _T_141 = 2'h0 == state2; // @[Conditional.scala 37:30]
  wire  _T_142 = io_dataReadBus_req_ready & io_dataReadBus_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_143 = 2'h1 == state2; // @[Conditional.scala 37:30]
  wire  _T_144 = 2'h2 == state2; // @[Conditional.scala 37:30]
  wire  _T_145 = io_mem_req_ready & io_mem_req_valid; // @[Decoupled.scala 40:37]
  wire  _T_147 = _T_145 | io_cohResp_valid; // @[Cache.scala 301:46]
  wire  _T_149 = _T_147 | hitReadBurst; // @[Cache.scala 301:67]
  wire [31:0] raddr = {io_in_bits_req_addr[31:3],3'h0}; // @[Cat.scala 29:58]
  wire [31:0] waddr = {meta_tag,addr_index,6'h0}; // @[Cat.scala 29:58]
  wire  _T_152 = state == 4'h1; // @[Cache.scala 309:23]
  wire  _T_153 = value_2 == 3'h7; // @[Cache.scala 310:29]
  wire [2:0] _T_154 = _T_153 ? 3'h7 : 3'h3; // @[Cache.scala 310:8]
  wire [2:0] cmd = _T_152 ? 3'h2 : _T_154; // @[Cache.scala 309:16]
  wire  _T_160 = state2 == 2'h2; // @[Cache.scala 316:89]
  wire  _T_161 = _T_118 & _T_160; // @[Cache.scala 316:78]
  reg  afterFirstRead; // @[Cache.scala 323:31]
  reg  alreadyOutFire; // @[Reg.scala 27:20]
  wire  _GEN_12 = io_out_valid | alreadyOutFire; // @[Reg.scala 28:19]
  wire  _T_165 = ~afterFirstRead; // @[Cache.scala 325:22]
  wire  _T_166 = io_mem_resp_ready & io_mem_resp_valid; // @[Decoupled.scala 40:37]
  wire  _T_167 = _T_165 & _T_166; // @[Cache.scala 325:38]
  wire  _T_168 = state == 4'h2; // @[Cache.scala 325:70]
  wire  readingFirst = _T_167 & _T_168; // @[Cache.scala 325:60]
  wire  _T_170 = state == 4'h6; // @[Cache.scala 327:52]
  wire  _T_171 = mmio ? _T_170 : readingFirst; // @[Cache.scala 327:39]
  reg [63:0] inRdataRegDemand; // @[Reg.scala 15:16]
  wire  _T_172 = state == 4'h0; // @[Cache.scala 330:31]
  wire  _T_173 = _T_172 & probe; // @[Cache.scala 330:43]
  wire  _T_176 = _T_119 & _T_160; // @[Cache.scala 331:46]
  wire  _T_180 = _T_119 & io_cohResp_valid; // @[Cache.scala 333:49]
  reg [2:0] _T_181; // @[Counter.scala 29:33]
  wire  _T_182 = _T_181 == 3'h7; // @[Counter.scala 38:24]
  wire [2:0] _T_184 = _T_181 + 3'h1; // @[Counter.scala 39:22]
  wire  releaseLast = _T_180 & _T_182; // @[Counter.scala 67:17]
  wire  respToL1Fire = hitReadBurst & _T_160; // @[Cache.scala 337:51]
  wire  _T_195 = _T_172 | _T_176; // @[Cache.scala 338:48]
  wire  _T_196 = _T_195 & hitReadBurst; // @[Cache.scala 338:96]
  reg [2:0] _T_198; // @[Counter.scala 29:33]
  wire  _T_199 = _T_198 == 3'h7; // @[Counter.scala 38:24]
  wire [2:0] _T_201 = _T_198 + 3'h1; // @[Counter.scala 39:22]
  wire  respToL1Last = _T_196 & _T_199; // @[Counter.scala 67:17]
  wire  _T_202 = 4'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_206 = addr_wordIndex == 3'h7; // @[Cache.scala 352:49]
  wire [2:0] _T_208 = addr_wordIndex + 3'h1; // @[Cache.scala 352:93]
  wire  _T_210 = miss | mmio; // @[Cache.scala 353:26]
  wire  _T_217 = 4'h5 == state; // @[Conditional.scala 37:30]
  wire  _T_219 = 4'h6 == state; // @[Conditional.scala 37:30]
  wire  _T_221 = 4'h8 == state; // @[Conditional.scala 37:30]
  wire  _T_223 = io_cohResp_valid | respToL1Fire; // @[Cache.scala 362:31]
  wire [2:0] _T_226 = value_1 + 3'h1; // @[Counter.scala 39:22]
  wire  _T_228 = probe & io_cohResp_valid; // @[Cache.scala 363:19]
  wire  _T_229 = _T_228 & releaseLast; // @[Cache.scala 363:40]
  wire  _T_230 = respToL1Fire & respToL1Last; // @[Cache.scala 363:71]
  wire  _T_231 = _T_229 | _T_230; // @[Cache.scala 363:55]
  wire  _T_232 = 4'h1 == state; // @[Conditional.scala 37:30]
  wire  _T_234 = 4'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_240 = io_mem_resp_bits_cmd == 4'h6; // @[SimpleBus.scala 91:26]
  wire  _GEN_33 = _T_166 | afterFirstRead; // @[Cache.scala 372:33]
  wire  _T_241 = 4'h3 == state; // @[Conditional.scala 37:30]
  wire [2:0] _T_245 = value_2 + 3'h1; // @[Counter.scala 39:22]
  wire  _T_246 = io_mem_req_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_248 = _T_246 & _T_145; // @[Cache.scala 382:43]
  wire  _T_249 = 4'h4 == state; // @[Conditional.scala 37:30]
  wire  _T_251 = 4'h7 == state; // @[Conditional.scala 37:30]
  wire [63:0] _T_255 = readingFirst ? wordMask : 64'h0; // @[Cache.scala 389:67]
  wire [63:0] _T_256 = io_in_bits_req_wdata & _T_255; // @[BitUtils.scala 32:13]
  wire [63:0] _T_257 = ~_T_255; // @[BitUtils.scala 32:38]
  wire [63:0] _T_258 = io_mem_resp_bits_rdata & _T_257; // @[BitUtils.scala 32:36]
  wire [63:0] dataRefill = _T_256 | _T_258; // @[BitUtils.scala 32:25]
  wire  dataRefillWriteBus_req_valid = _T_168 & _T_166; // @[Cache.scala 391:39]
  wire  metaRefillWriteBus_req_valid = dataRefillWriteBus_req_valid & _T_240; // @[Cache.scala 399:61]
  wire  _T_283 = dataRefillWriteBus_req_valid & _T_8; // @[Cache.scala 409:59]
  wire [2:0] _T_285 = _T_240 ? 3'h6 : 3'h2; // @[Cache.scala 412:29]
  wire  _T_288 = _T_88 | _T_87; // @[Cache.scala 413:35]
  wire [63:0] _T_289 = hit ? dataRead : inRdataRegDemand; // @[Cache.scala 415:31]
  wire  _T_291 = hitReadBurst & _T_119; // @[Cache.scala 417:30]
  wire [2:0] _T_292 = respToL1Last ? 3'h6 : 3'h2; // @[Cache.scala 420:29]
  wire [63:0] _GEN_76 = _T_291 ? _T_137 : _T_289; // @[Cache.scala 417:54]
  wire [3:0] _GEN_77 = _T_291 ? {{1'd0}, _T_292} : io_in_bits_req_cmd; // @[Cache.scala 417:54]
  wire [63:0] _GEN_78 = _T_288 ? _T_289 : _GEN_76; // @[Cache.scala 413:75]
  wire  _T_297 = ~hit; // @[Cache.scala 433:34]
  wire  _T_298 = state == 4'h7; // @[Cache.scala 433:48]
  wire  _T_299 = _T_297 & _T_298; // @[Cache.scala 433:39]
  wire  _T_300 = hit | _T_299; // @[Cache.scala 433:31]
  wire  _T_301 = io_in_bits_req_cmd[0] & _T_300; // @[Cache.scala 433:23]
  wire  _T_307 = _T_301 | _T_283; // @[Cache.scala 433:8]
  wire  _T_310 = _T_230 & _T_119; // @[Cache.scala 433:194]
  wire  _T_311 = _T_307 | _T_310; // @[Cache.scala 433:161]
  wire  _T_313 = io_in_bits_req_cmd[0] | mmio; // @[Cache.scala 434:60]
  wire  _T_315 = ~alreadyOutFire; // @[Cache.scala 434:110]
  wire  _T_316 = afterFirstRead & _T_315; // @[Cache.scala 434:107]
  wire  _T_317 = _T_313 ? _T_298 : _T_316; // @[Cache.scala 434:45]
  wire  _T_318 = hit | _T_317; // @[Cache.scala 434:28]
  wire  _T_319 = probe ? 1'h0 : _T_318; // @[Cache.scala 434:8]
  wire  _T_320 = io_in_bits_req_cmd[1] ? _T_311 : _T_319; // @[Cache.scala 432:37]
  wire  _T_325 = _T_119 & releaseLast; // @[Cache.scala 441:100]
  wire  _T_326 = miss ? _T_172 : _T_325; // @[Cache.scala 441:53]
  wire  _T_327 = io_cohResp_valid & _T_326; // @[Cache.scala 441:47]
  wire  _T_329 = hit | io_in_bits_req_cmd[0]; // @[Cache.scala 442:13]
  wire  _T_334 = _T_298 & _GEN_12; // @[Cache.scala 442:70]
  wire  _T_335 = _T_329 ? io_out_valid : _T_334; // @[Cache.scala 442:8]
  wire  _T_338 = ~hitReadBurst; // @[Cache.scala 445:55]
  wire  _T_339 = _T_172 & _T_338; // @[Cache.scala 445:52]
  wire  _T_341 = ~miss; // @[Cache.scala 445:73]
  wire  _T_342 = _T_339 & _T_341; // @[Cache.scala 445:70]
  wire  _T_343 = ~probe; // @[Cache.scala 445:82]
  wire  _T_352 = metaHitWriteBus_req_valid & metaRefillWriteBus_req_valid; // @[Cache.scala 448:38]
  wire  _T_353 = ~_T_352; // @[Cache.scala 448:10]
  wire  _T_355 = _T_353 | reset; // @[Cache.scala 448:9]
  wire  _T_356 = ~_T_355; // @[Cache.scala 448:9]
  wire  _T_357 = hitWrite & dataRefillWriteBus_req_valid; // @[Cache.scala 449:38]
  wire  _T_358 = ~_T_357; // @[Cache.scala 449:10]
  wire  _T_360 = _T_358 | reset; // @[Cache.scala 449:9]
  wire  _T_361 = ~_T_360; // @[Cache.scala 449:9]
  Arbiter_10 metaWriteArb ( // @[Cache.scala 241:28]
    .io_in_0_valid(metaWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(metaWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_tag(metaWriteArb_io_in_0_bits_data_tag),
    .io_in_0_bits_waymask(metaWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(metaWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(metaWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_tag(metaWriteArb_io_in_1_bits_data_tag),
    .io_in_1_bits_data_dirty(metaWriteArb_io_in_1_bits_data_dirty),
    .io_in_1_bits_waymask(metaWriteArb_io_in_1_bits_waymask),
    .io_out_valid(metaWriteArb_io_out_valid),
    .io_out_bits_setIdx(metaWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_tag(metaWriteArb_io_out_bits_data_tag),
    .io_out_bits_data_dirty(metaWriteArb_io_out_bits_data_dirty),
    .io_out_bits_waymask(metaWriteArb_io_out_bits_waymask)
  );
  Arbiter_11 dataWriteArb ( // @[Cache.scala 242:28]
    .io_in_0_valid(dataWriteArb_io_in_0_valid),
    .io_in_0_bits_setIdx(dataWriteArb_io_in_0_bits_setIdx),
    .io_in_0_bits_data_data(dataWriteArb_io_in_0_bits_data_data),
    .io_in_0_bits_waymask(dataWriteArb_io_in_0_bits_waymask),
    .io_in_1_valid(dataWriteArb_io_in_1_valid),
    .io_in_1_bits_setIdx(dataWriteArb_io_in_1_bits_setIdx),
    .io_in_1_bits_data_data(dataWriteArb_io_in_1_bits_data_data),
    .io_in_1_bits_waymask(dataWriteArb_io_in_1_bits_waymask),
    .io_out_valid(dataWriteArb_io_out_valid),
    .io_out_bits_setIdx(dataWriteArb_io_out_bits_setIdx),
    .io_out_bits_data_data(dataWriteArb_io_out_bits_data_data),
    .io_out_bits_waymask(dataWriteArb_io_out_bits_waymask)
  );
  assign io_in_ready = _T_342 & _T_343; // @[Cache.scala 445:15]
  assign io_out_valid = io_in_valid & _T_320; // @[Cache.scala 432:16]
  assign io_out_bits_cmd = _T_283 ? {{1'd0}, _T_285} : _GEN_77; // @[Cache.scala 412:23 Cache.scala 420:23 Cache.scala 423:23]
  assign io_out_bits_rdata = _T_283 ? dataRefill : _GEN_78; // @[Cache.scala 411:25 Cache.scala 415:25 Cache.scala 419:25 Cache.scala 422:25]
  assign io_isFinish = probe ? _T_327 : _T_335; // @[Cache.scala 441:15]
  assign io_dataReadBus_req_valid = _T_120 & _T_121; // @[SRAMTemplate.scala 53:20]
  assign io_dataReadBus_req_bits_setIdx = {addr_index,_T_124}; // @[SRAMTemplate.scala 26:17]
  assign io_dataWriteBus_req_valid = dataWriteArb_io_out_valid; // @[Cache.scala 396:23]
  assign io_dataWriteBus_req_bits_setIdx = dataWriteArb_io_out_bits_setIdx; // @[Cache.scala 396:23]
  assign io_dataWriteBus_req_bits_data_data = dataWriteArb_io_out_bits_data_data; // @[Cache.scala 396:23]
  assign io_dataWriteBus_req_bits_waymask = dataWriteArb_io_out_bits_waymask; // @[Cache.scala 396:23]
  assign io_metaWriteBus_req_valid = metaWriteArb_io_out_valid; // @[Cache.scala 406:23]
  assign io_metaWriteBus_req_bits_setIdx = metaWriteArb_io_out_bits_setIdx; // @[Cache.scala 406:23]
  assign io_metaWriteBus_req_bits_data_tag = metaWriteArb_io_out_bits_data_tag; // @[Cache.scala 406:23]
  assign io_metaWriteBus_req_bits_data_dirty = metaWriteArb_io_out_bits_data_dirty; // @[Cache.scala 406:23]
  assign io_metaWriteBus_req_bits_waymask = metaWriteArb_io_out_bits_waymask; // @[Cache.scala 406:23]
  assign io_mem_req_valid = _T_152 | _T_161; // @[Cache.scala 316:20]
  assign io_mem_req_bits_addr = _T_152 ? raddr : waddr; // @[SimpleBus.scala 64:15]
  assign io_mem_req_bits_cmd = {{1'd0}, cmd}; // @[SimpleBus.scala 65:14]
  assign io_mem_req_bits_wdata = _T_136 | _T_134; // @[SimpleBus.scala 67:16]
  assign io_mem_resp_ready = 1'h1; // @[Cache.scala 315:21]
  assign io_cohResp_valid = _T_173 | _T_176; // @[Cache.scala 330:20]
  assign io_dataReadRespToL1 = hitReadBurst & _T_195; // @[Cache.scala 446:23]
  assign metaWriteArb_io_in_0_valid = hitWrite & _T_105; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_0_bits_setIdx = io_in_bits_req_addr[14:6]; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_0_bits_data_tag = _T_27[18:2]; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 404:25]
  assign metaWriteArb_io_in_1_valid = dataRefillWriteBus_req_valid & _T_240; // @[Cache.scala 405:25]
  assign metaWriteArb_io_in_1_bits_setIdx = io_in_bits_req_addr[14:6]; // @[Cache.scala 405:25]
  assign metaWriteArb_io_in_1_bits_data_tag = io_in_bits_req_addr[31:15]; // @[Cache.scala 405:25]
  assign metaWriteArb_io_in_1_bits_data_dirty = io_in_bits_req_cmd[0]; // @[Cache.scala 405:25]
  assign metaWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 405:25]
  assign dataWriteArb_io_in_0_valid = hit & io_in_bits_req_cmd[0]; // @[Cache.scala 394:25]
  assign dataWriteArb_io_in_0_bits_setIdx = {addr_index,_T_103}; // @[Cache.scala 394:25]
  assign dataWriteArb_io_in_0_bits_data_data = _T_96 | _T_98; // @[Cache.scala 394:25]
  assign dataWriteArb_io_in_0_bits_waymask = io_in_bits_waymask; // @[Cache.scala 394:25]
  assign dataWriteArb_io_in_1_valid = _T_168 & _T_166; // @[Cache.scala 395:25]
  assign dataWriteArb_io_in_1_bits_setIdx = {addr_index,value_1}; // @[Cache.scala 395:25]
  assign dataWriteArb_io_in_1_bits_data_data = _T_256 | _T_258; // @[Cache.scala 395:25]
  assign dataWriteArb_io_in_1_bits_waymask = io_in_bits_waymask; // @[Cache.scala 395:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  value = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  state = _RAND_1[3:0];
  _RAND_2 = {1{`RANDOM}};
  value_1 = _RAND_2[2:0];
  _RAND_3 = {1{`RANDOM}};
  value_2 = _RAND_3[2:0];
  _RAND_4 = {1{`RANDOM}};
  state2 = _RAND_4[1:0];
  _RAND_5 = {2{`RANDOM}};
  dataWay_0_data = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  dataWay_1_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  dataWay_2_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  dataWay_3_data = _RAND_8[63:0];
  _RAND_9 = {1{`RANDOM}};
  afterFirstRead = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  alreadyOutFire = _RAND_10[0:0];
  _RAND_11 = {2{`RANDOM}};
  inRdataRegDemand = _RAND_11[63:0];
  _RAND_12 = {1{`RANDOM}};
  _T_181 = _RAND_12[2:0];
  _RAND_13 = {1{`RANDOM}};
  _T_198 = _RAND_13[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      value <= 3'h0;
    end else if (_T_202) begin
      if (_T_90) begin
        value <= _T_93;
      end
    end else if (_T_217) begin
      if (_T_90) begin
        value <= _T_93;
      end
    end else if (_T_219) begin
      if (_T_90) begin
        value <= _T_93;
      end
    end else if (_T_221) begin
      if (_T_90) begin
        value <= _T_93;
      end
    end else if (_T_232) begin
      value <= _GEN_0;
    end else if (_T_234) begin
      if (_T_166) begin
        if (_T_87) begin
          value <= 3'h0;
        end else begin
          value <= _GEN_0;
        end
      end else begin
        value <= _GEN_0;
      end
    end else begin
      value <= _GEN_0;
    end
    if (reset) begin
      state <= 4'h0;
    end else if (_T_202) begin
      if (probe) begin
        if (io_cohResp_valid) begin
          if (hit) begin
            state <= 4'h8;
          end else begin
            state <= 4'h0;
          end
        end
      end else if (hitReadBurst) begin
        state <= 4'h8;
      end else if (_T_210) begin
        if (mmio) begin
          state <= 4'h5;
        end else if (meta_dirty) begin
          state <= 4'h3;
        end else begin
          state <= 4'h1;
        end
      end
    end else if (!(_T_217)) begin
      if (!(_T_219)) begin
        if (_T_221) begin
          if (_T_231) begin
            state <= 4'h0;
          end
        end else if (_T_232) begin
          if (_T_145) begin
            state <= 4'h2;
          end
        end else if (_T_234) begin
          if (_T_166) begin
            if (_T_240) begin
              state <= 4'h7;
            end
          end
        end else if (_T_241) begin
          if (_T_248) begin
            state <= 4'h4;
          end
        end else if (_T_249) begin
          if (_T_166) begin
            state <= 4'h1;
          end
        end else if (_T_251) begin
          if (_GEN_12) begin
            state <= 4'h0;
          end
        end
      end
    end
    if (reset) begin
      value_1 <= 3'h0;
    end else if (_T_202) begin
      if (probe) begin
        if (io_cohResp_valid) begin
          value_1 <= addr_wordIndex;
        end
      end else if (hitReadBurst) begin
        if (_T_206) begin
          value_1 <= 3'h0;
        end else begin
          value_1 <= _T_208;
        end
      end
    end else if (!(_T_217)) begin
      if (!(_T_219)) begin
        if (_T_221) begin
          if (_T_223) begin
            value_1 <= _T_226;
          end
        end else if (_T_232) begin
          if (_T_145) begin
            value_1 <= addr_wordIndex;
          end
        end else if (_T_234) begin
          if (_T_166) begin
            value_1 <= _T_226;
          end
        end
      end
    end
    if (reset) begin
      value_2 <= 3'h0;
    end else if (!(_T_202)) begin
      if (!(_T_217)) begin
        if (!(_T_219)) begin
          if (!(_T_221)) begin
            if (!(_T_232)) begin
              if (!(_T_234)) begin
                if (_T_241) begin
                  if (_T_145) begin
                    value_2 <= _T_245;
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      state2 <= 2'h0;
    end else if (_T_141) begin
      if (_T_142) begin
        state2 <= 2'h1;
      end
    end else if (_T_143) begin
      state2 <= 2'h2;
    end else if (_T_144) begin
      if (_T_149) begin
        state2 <= 2'h0;
      end
    end
    if (_T_126) begin
      dataWay_0_data <= io_dataReadBus_resp_data_0_data;
    end
    if (_T_126) begin
      dataWay_1_data <= io_dataReadBus_resp_data_1_data;
    end
    if (_T_126) begin
      dataWay_2_data <= io_dataReadBus_resp_data_2_data;
    end
    if (_T_126) begin
      dataWay_3_data <= io_dataReadBus_resp_data_3_data;
    end
    if (reset) begin
      afterFirstRead <= 1'h0;
    end else if (_T_202) begin
      afterFirstRead <= 1'h0;
    end else if (!(_T_217)) begin
      if (!(_T_219)) begin
        if (!(_T_221)) begin
          if (!(_T_232)) begin
            if (_T_234) begin
              afterFirstRead <= _GEN_33;
            end
          end
        end
      end
    end
    if (reset) begin
      alreadyOutFire <= 1'h0;
    end else if (_T_202) begin
      alreadyOutFire <= 1'h0;
    end else begin
      alreadyOutFire <= _GEN_12;
    end
    if (_T_171) begin
      if (mmio) begin
        inRdataRegDemand <= 64'h0;
      end else begin
        inRdataRegDemand <= io_mem_resp_bits_rdata;
      end
    end
    if (reset) begin
      _T_181 <= 3'h0;
    end else if (_T_180) begin
      _T_181 <= _T_184;
    end
    if (reset) begin
      _T_198 <= 3'h0;
    end else if (_T_196) begin
      _T_198 <= _T_201;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_36) begin
          $fwrite(32'h80000002,"Assertion failed: MMIO request should not hit in cache\n    at Cache.scala:252 assert(!(mmio && hit), \"MMIO request should not hit in cache\")\n"); // @[Cache.scala 252:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_36) begin
          $fatal; // @[Cache.scala 252:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_356) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Cache.scala:448 assert(!(metaHitWriteBus.req.valid && metaRefillWriteBus.req.valid))\n"); // @[Cache.scala 448:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_356) begin
          $fatal; // @[Cache.scala 448:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_361) begin
          $fwrite(32'h80000002,"Assertion failed\n    at Cache.scala:449 assert(!(dataHitWriteBus.req.valid && dataRefillWriteBus.req.valid))\n"); // @[Cache.scala 449:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_361) begin
          $fatal; // @[Cache.scala 449:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module SRAMTemplate_5(
  input         clock,
  input         reset,
  output        io_rreq_ready,
  input         io_rreq_valid,
  input  [8:0]  io_rreq_bits_setIdx,
  output [16:0] io_rresp_data_0_tag,
  output        io_rresp_data_0_valid,
  output        io_rresp_data_0_dirty,
  output [16:0] io_rresp_data_1_tag,
  output        io_rresp_data_1_valid,
  output        io_rresp_data_1_dirty,
  output [16:0] io_rresp_data_2_tag,
  output        io_rresp_data_2_valid,
  output        io_rresp_data_2_dirty,
  output [16:0] io_rresp_data_3_tag,
  output        io_rresp_data_3_valid,
  output        io_rresp_data_3_dirty,
  input         io_wreq_valid,
  input  [8:0]  io_wreq_bits_setIdx,
  input  [16:0] io_wreq_bits_data_tag,
  input         io_wreq_bits_data_dirty,
  input  [3:0]  io_wreq_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire [8:0] array_RW0_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_en; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_clk; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmode; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_RW0_wdata_0; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_RW0_wdata_1; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_RW0_wdata_2; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_RW0_wdata_3; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_RW0_rdata_0; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_RW0_rdata_1; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_RW0_rdata_2; // @[SRAMTemplate.scala 76:26]
  wire [18:0] array_RW0_rdata_3; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_0; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_1; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_2; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_3; // @[SRAMTemplate.scala 76:26]
  reg  resetState; // @[SRAMTemplate.scala 80:30]
  reg [8:0] resetSet; // @[Counter.scala 29:33]
  wire  _T_3 = resetSet == 9'h1ff; // @[Counter.scala 38:24]
  wire [8:0] _T_5 = resetSet + 9'h1; // @[Counter.scala 39:22]
  wire  _GEN_1 = resetState & _T_3; // @[Counter.scala 67:17]
  wire  _GEN_2 = _GEN_1 ? 1'h0 : resetState; // @[SRAMTemplate.scala 82:24]
  wire  wen = io_wreq_valid | resetState; // @[SRAMTemplate.scala 88:52]
  wire  _T_6 = ~wen; // @[SRAMTemplate.scala 89:41]
  wire  realRen = io_rreq_valid & _T_6; // @[SRAMTemplate.scala 89:38]
  wire [8:0] setIdx = resetState ? resetSet : io_wreq_bits_setIdx; // @[SRAMTemplate.scala 91:19]
  wire [18:0] _T_9 = {io_wreq_bits_data_tag,1'h1,io_wreq_bits_data_dirty}; // @[SRAMTemplate.scala 92:78]
  wire [3:0] waymask = resetState ? 4'hf : io_wreq_bits_waymask; // @[SRAMTemplate.scala 93:20]
  wire [18:0] _T_22 = array_RW0_rdata_0;
  wire [18:0] _T_26 = array_RW0_rdata_1;
  wire [18:0] _T_30 = array_RW0_rdata_2;
  wire [18:0] _T_34 = array_RW0_rdata_3;
  wire  _T_39 = ~resetState; // @[SRAMTemplate.scala 101:21]
  array_2 array ( // @[SRAMTemplate.scala 76:26]
    .RW0_addr(array_RW0_addr),
    .RW0_en(array_RW0_en),
    .RW0_clk(array_RW0_clk),
    .RW0_wmode(array_RW0_wmode),
    .RW0_wdata_0(array_RW0_wdata_0),
    .RW0_wdata_1(array_RW0_wdata_1),
    .RW0_wdata_2(array_RW0_wdata_2),
    .RW0_wdata_3(array_RW0_wdata_3),
    .RW0_rdata_0(array_RW0_rdata_0),
    .RW0_rdata_1(array_RW0_rdata_1),
    .RW0_rdata_2(array_RW0_rdata_2),
    .RW0_rdata_3(array_RW0_rdata_3),
    .RW0_wmask_0(array_RW0_wmask_0),
    .RW0_wmask_1(array_RW0_wmask_1),
    .RW0_wmask_2(array_RW0_wmask_2),
    .RW0_wmask_3(array_RW0_wmask_3)
  );
  assign io_rreq_ready = _T_39 & _T_6; // @[SRAMTemplate.scala 101:18]
  assign io_rresp_data_0_tag = _T_22[18:2]; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_0_valid = _T_22[1]; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_0_dirty = _T_22[0]; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_1_tag = _T_26[18:2]; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_1_valid = _T_26[1]; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_1_dirty = _T_26[0]; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_2_tag = _T_30[18:2]; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_2_valid = _T_30[1]; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_2_dirty = _T_30[0]; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_3_tag = _T_34[18:2]; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_3_valid = _T_34[1]; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_3_dirty = _T_34[0]; // @[SRAMTemplate.scala 99:18]
  assign array_RW0_wdata_0 = resetState ? 19'h0 : _T_9;
  assign array_RW0_wdata_1 = resetState ? 19'h0 : _T_9;
  assign array_RW0_wdata_2 = resetState ? 19'h0 : _T_9;
  assign array_RW0_wdata_3 = resetState ? 19'h0 : _T_9;
  assign array_RW0_wmask_0 = waymask[0];
  assign array_RW0_wmask_1 = waymask[1];
  assign array_RW0_wmask_2 = waymask[2];
  assign array_RW0_wmask_3 = waymask[3];
  assign array_RW0_wmode = io_wreq_valid | resetState;
  assign array_RW0_clk = clock;
  assign array_RW0_en = realRen | wen;
  assign array_RW0_addr = wen ? setIdx : io_rreq_bits_setIdx;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  resetState = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  resetSet = _RAND_1[8:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    resetState <= reset | _GEN_2;
    if (reset) begin
      resetSet <= 9'h0;
    end else if (resetState) begin
      resetSet <= _T_5;
    end
  end
endmodule
module Arbiter_12(
  output       io_in_0_ready,
  input        io_in_0_valid,
  input  [8:0] io_in_0_bits_setIdx,
  input        io_out_ready,
  output       io_out_valid,
  output [8:0] io_out_bits_setIdx
);
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = io_in_0_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_setIdx = io_in_0_bits_setIdx; // @[Arbiter.scala 124:15]
endmodule
module SRAMTemplateWithArbiter_4(
  input         clock,
  input         reset,
  output        io_r0_req_ready,
  input         io_r0_req_valid,
  input  [8:0]  io_r0_req_bits_setIdx,
  output [16:0] io_r0_resp_data_0_tag,
  output        io_r0_resp_data_0_valid,
  output        io_r0_resp_data_0_dirty,
  output [16:0] io_r0_resp_data_1_tag,
  output        io_r0_resp_data_1_valid,
  output        io_r0_resp_data_1_dirty,
  output [16:0] io_r0_resp_data_2_tag,
  output        io_r0_resp_data_2_valid,
  output        io_r0_resp_data_2_dirty,
  output [16:0] io_r0_resp_data_3_tag,
  output        io_r0_resp_data_3_valid,
  output        io_r0_resp_data_3_dirty,
  input         io_wreq_valid,
  input  [8:0]  io_wreq_bits_setIdx,
  input  [16:0] io_wreq_bits_data_tag,
  input         io_wreq_bits_data_dirty,
  input  [3:0]  io_wreq_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire  ram_clock; // @[SRAMTemplate.scala 121:19]
  wire  ram_reset; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rreq_ready; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rreq_valid; // @[SRAMTemplate.scala 121:19]
  wire [8:0] ram_io_rreq_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [16:0] ram_io_rresp_data_0_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_0_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_0_dirty; // @[SRAMTemplate.scala 121:19]
  wire [16:0] ram_io_rresp_data_1_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_1_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_1_dirty; // @[SRAMTemplate.scala 121:19]
  wire [16:0] ram_io_rresp_data_2_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_2_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_2_dirty; // @[SRAMTemplate.scala 121:19]
  wire [16:0] ram_io_rresp_data_3_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_3_valid; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rresp_data_3_dirty; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_wreq_valid; // @[SRAMTemplate.scala 121:19]
  wire [8:0] ram_io_wreq_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [16:0] ram_io_wreq_bits_data_tag; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_wreq_bits_data_dirty; // @[SRAMTemplate.scala 121:19]
  wire [3:0] ram_io_wreq_bits_waymask; // @[SRAMTemplate.scala 121:19]
  wire  readArb_io_in_0_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_0_valid; // @[SRAMTemplate.scala 124:23]
  wire [8:0] readArb_io_in_0_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_valid; // @[SRAMTemplate.scala 124:23]
  wire [8:0] readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  reg  _T_1; // @[SRAMTemplate.scala 130:58]
  reg [16:0] _T_3_0_tag; // @[Reg.scala 27:20]
  reg  _T_3_0_valid; // @[Reg.scala 27:20]
  reg  _T_3_0_dirty; // @[Reg.scala 27:20]
  reg [16:0] _T_3_1_tag; // @[Reg.scala 27:20]
  reg  _T_3_1_valid; // @[Reg.scala 27:20]
  reg  _T_3_1_dirty; // @[Reg.scala 27:20]
  reg [16:0] _T_3_2_tag; // @[Reg.scala 27:20]
  reg  _T_3_2_valid; // @[Reg.scala 27:20]
  reg  _T_3_2_dirty; // @[Reg.scala 27:20]
  reg [16:0] _T_3_3_tag; // @[Reg.scala 27:20]
  reg  _T_3_3_valid; // @[Reg.scala 27:20]
  reg  _T_3_3_dirty; // @[Reg.scala 27:20]
  SRAMTemplate_5 ram ( // @[SRAMTemplate.scala 121:19]
    .clock(ram_clock),
    .reset(ram_reset),
    .io_rreq_ready(ram_io_rreq_ready),
    .io_rreq_valid(ram_io_rreq_valid),
    .io_rreq_bits_setIdx(ram_io_rreq_bits_setIdx),
    .io_rresp_data_0_tag(ram_io_rresp_data_0_tag),
    .io_rresp_data_0_valid(ram_io_rresp_data_0_valid),
    .io_rresp_data_0_dirty(ram_io_rresp_data_0_dirty),
    .io_rresp_data_1_tag(ram_io_rresp_data_1_tag),
    .io_rresp_data_1_valid(ram_io_rresp_data_1_valid),
    .io_rresp_data_1_dirty(ram_io_rresp_data_1_dirty),
    .io_rresp_data_2_tag(ram_io_rresp_data_2_tag),
    .io_rresp_data_2_valid(ram_io_rresp_data_2_valid),
    .io_rresp_data_2_dirty(ram_io_rresp_data_2_dirty),
    .io_rresp_data_3_tag(ram_io_rresp_data_3_tag),
    .io_rresp_data_3_valid(ram_io_rresp_data_3_valid),
    .io_rresp_data_3_dirty(ram_io_rresp_data_3_dirty),
    .io_wreq_valid(ram_io_wreq_valid),
    .io_wreq_bits_setIdx(ram_io_wreq_bits_setIdx),
    .io_wreq_bits_data_tag(ram_io_wreq_bits_data_tag),
    .io_wreq_bits_data_dirty(ram_io_wreq_bits_data_dirty),
    .io_wreq_bits_waymask(ram_io_wreq_bits_waymask)
  );
  Arbiter_12 readArb ( // @[SRAMTemplate.scala 124:23]
    .io_in_0_ready(readArb_io_in_0_ready),
    .io_in_0_valid(readArb_io_in_0_valid),
    .io_in_0_bits_setIdx(readArb_io_in_0_bits_setIdx),
    .io_out_ready(readArb_io_out_ready),
    .io_out_valid(readArb_io_out_valid),
    .io_out_bits_setIdx(readArb_io_out_bits_setIdx)
  );
  assign io_r0_req_ready = readArb_io_in_0_ready; // @[SRAMTemplate.scala 125:17]
  assign io_r0_resp_data_0_tag = _T_1 ? ram_io_rresp_data_0_tag : _T_3_0_tag; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_0_valid = _T_1 ? ram_io_rresp_data_0_valid : _T_3_0_valid; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_0_dirty = _T_1 ? ram_io_rresp_data_0_dirty : _T_3_0_dirty; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_1_tag = _T_1 ? ram_io_rresp_data_1_tag : _T_3_1_tag; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_1_valid = _T_1 ? ram_io_rresp_data_1_valid : _T_3_1_valid; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_1_dirty = _T_1 ? ram_io_rresp_data_1_dirty : _T_3_1_dirty; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_2_tag = _T_1 ? ram_io_rresp_data_2_tag : _T_3_2_tag; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_2_valid = _T_1 ? ram_io_rresp_data_2_valid : _T_3_2_valid; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_2_dirty = _T_1 ? ram_io_rresp_data_2_dirty : _T_3_2_dirty; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_3_tag = _T_1 ? ram_io_rresp_data_3_tag : _T_3_3_tag; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_3_valid = _T_1 ? ram_io_rresp_data_3_valid : _T_3_3_valid; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_3_dirty = _T_1 ? ram_io_rresp_data_3_dirty : _T_3_3_dirty; // @[SRAMTemplate.scala 130:17]
  assign ram_clock = clock;
  assign ram_reset = reset;
  assign ram_io_rreq_valid = readArb_io_out_valid; // @[SRAMTemplate.scala 126:16]
  assign ram_io_rreq_bits_setIdx = readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 126:16]
  assign ram_io_wreq_valid = io_wreq_valid; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_setIdx = io_wreq_bits_setIdx; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_data_tag = io_wreq_bits_data_tag; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_data_dirty = io_wreq_bits_data_dirty; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_waymask = io_wreq_bits_waymask; // @[SRAMTemplate.scala 122:12]
  assign readArb_io_in_0_valid = io_r0_req_valid; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_0_bits_setIdx = io_r0_req_bits_setIdx; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_out_ready = ram_io_rreq_ready; // @[SRAMTemplate.scala 126:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _T_3_0_tag = _RAND_1[16:0];
  _RAND_2 = {1{`RANDOM}};
  _T_3_0_valid = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  _T_3_0_dirty = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_3_1_tag = _RAND_4[16:0];
  _RAND_5 = {1{`RANDOM}};
  _T_3_1_valid = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_3_1_dirty = _RAND_6[0:0];
  _RAND_7 = {1{`RANDOM}};
  _T_3_2_tag = _RAND_7[16:0];
  _RAND_8 = {1{`RANDOM}};
  _T_3_2_valid = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  _T_3_2_dirty = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  _T_3_3_tag = _RAND_10[16:0];
  _RAND_11 = {1{`RANDOM}};
  _T_3_3_valid = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _T_3_3_dirty = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_1 <= io_r0_req_ready & io_r0_req_valid;
    if (reset) begin
      _T_3_0_tag <= 17'h0;
    end else if (_T_1) begin
      _T_3_0_tag <= ram_io_rresp_data_0_tag;
    end
    if (reset) begin
      _T_3_0_valid <= 1'h0;
    end else if (_T_1) begin
      _T_3_0_valid <= ram_io_rresp_data_0_valid;
    end
    if (reset) begin
      _T_3_0_dirty <= 1'h0;
    end else if (_T_1) begin
      _T_3_0_dirty <= ram_io_rresp_data_0_dirty;
    end
    if (reset) begin
      _T_3_1_tag <= 17'h0;
    end else if (_T_1) begin
      _T_3_1_tag <= ram_io_rresp_data_1_tag;
    end
    if (reset) begin
      _T_3_1_valid <= 1'h0;
    end else if (_T_1) begin
      _T_3_1_valid <= ram_io_rresp_data_1_valid;
    end
    if (reset) begin
      _T_3_1_dirty <= 1'h0;
    end else if (_T_1) begin
      _T_3_1_dirty <= ram_io_rresp_data_1_dirty;
    end
    if (reset) begin
      _T_3_2_tag <= 17'h0;
    end else if (_T_1) begin
      _T_3_2_tag <= ram_io_rresp_data_2_tag;
    end
    if (reset) begin
      _T_3_2_valid <= 1'h0;
    end else if (_T_1) begin
      _T_3_2_valid <= ram_io_rresp_data_2_valid;
    end
    if (reset) begin
      _T_3_2_dirty <= 1'h0;
    end else if (_T_1) begin
      _T_3_2_dirty <= ram_io_rresp_data_2_dirty;
    end
    if (reset) begin
      _T_3_3_tag <= 17'h0;
    end else if (_T_1) begin
      _T_3_3_tag <= ram_io_rresp_data_3_tag;
    end
    if (reset) begin
      _T_3_3_valid <= 1'h0;
    end else if (_T_1) begin
      _T_3_3_valid <= ram_io_rresp_data_3_valid;
    end
    if (reset) begin
      _T_3_3_dirty <= 1'h0;
    end else if (_T_1) begin
      _T_3_3_dirty <= ram_io_rresp_data_3_dirty;
    end
  end
endmodule
module SRAMTemplate_6(
  input         clock,
  output        io_rreq_ready,
  input         io_rreq_valid,
  input  [11:0] io_rreq_bits_setIdx,
  output [63:0] io_rresp_data_0_data,
  output [63:0] io_rresp_data_1_data,
  output [63:0] io_rresp_data_2_data,
  output [63:0] io_rresp_data_3_data,
  input         io_wreq_valid,
  input  [11:0] io_wreq_bits_setIdx,
  input  [63:0] io_wreq_bits_data_data,
  input  [3:0]  io_wreq_bits_waymask
);
  wire [11:0] array_RW0_addr; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_en; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_clk; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmode; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_wdata_0; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_wdata_1; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_wdata_2; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_wdata_3; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_rdata_0; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_rdata_1; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_rdata_2; // @[SRAMTemplate.scala 76:26]
  wire [63:0] array_RW0_rdata_3; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_0; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_1; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_2; // @[SRAMTemplate.scala 76:26]
  wire  array_RW0_wmask_3; // @[SRAMTemplate.scala 76:26]
  wire  _T = ~io_wreq_valid; // @[SRAMTemplate.scala 89:41]
  wire  realRen = io_rreq_valid & _T; // @[SRAMTemplate.scala 89:38]
  array_3 array ( // @[SRAMTemplate.scala 76:26]
    .RW0_addr(array_RW0_addr),
    .RW0_en(array_RW0_en),
    .RW0_clk(array_RW0_clk),
    .RW0_wmode(array_RW0_wmode),
    .RW0_wdata_0(array_RW0_wdata_0),
    .RW0_wdata_1(array_RW0_wdata_1),
    .RW0_wdata_2(array_RW0_wdata_2),
    .RW0_wdata_3(array_RW0_wdata_3),
    .RW0_rdata_0(array_RW0_rdata_0),
    .RW0_rdata_1(array_RW0_rdata_1),
    .RW0_rdata_2(array_RW0_rdata_2),
    .RW0_rdata_3(array_RW0_rdata_3),
    .RW0_wmask_0(array_RW0_wmask_0),
    .RW0_wmask_1(array_RW0_wmask_1),
    .RW0_wmask_2(array_RW0_wmask_2),
    .RW0_wmask_3(array_RW0_wmask_3)
  );
  assign io_rreq_ready = ~io_wreq_valid; // @[SRAMTemplate.scala 101:18]
  assign io_rresp_data_0_data = array_RW0_rdata_0; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_1_data = array_RW0_rdata_1; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_2_data = array_RW0_rdata_2; // @[SRAMTemplate.scala 99:18]
  assign io_rresp_data_3_data = array_RW0_rdata_3; // @[SRAMTemplate.scala 99:18]
  assign array_RW0_wdata_0 = io_wreq_bits_data_data;
  assign array_RW0_wdata_1 = io_wreq_bits_data_data;
  assign array_RW0_wdata_2 = io_wreq_bits_data_data;
  assign array_RW0_wdata_3 = io_wreq_bits_data_data;
  assign array_RW0_wmask_0 = io_wreq_bits_waymask[0];
  assign array_RW0_wmask_1 = io_wreq_bits_waymask[1];
  assign array_RW0_wmask_2 = io_wreq_bits_waymask[2];
  assign array_RW0_wmask_3 = io_wreq_bits_waymask[3];
  assign array_RW0_wmode = io_wreq_valid;
  assign array_RW0_clk = clock;
  assign array_RW0_en = realRen | io_wreq_valid;
  assign array_RW0_addr = io_wreq_valid ? io_wreq_bits_setIdx : io_rreq_bits_setIdx;
endmodule
module Arbiter_13(
  output        io_in_0_ready,
  input         io_in_0_valid,
  input  [11:0] io_in_0_bits_setIdx,
  output        io_in_1_ready,
  input         io_in_1_valid,
  input  [11:0] io_in_1_bits_setIdx,
  input         io_out_ready,
  output        io_out_valid,
  output [11:0] io_out_bits_setIdx
);
  wire  grant_1 = ~io_in_0_valid; // @[Arbiter.scala 31:78]
  wire  _T_2 = ~grant_1; // @[Arbiter.scala 135:19]
  assign io_in_0_ready = io_out_ready; // @[Arbiter.scala 134:14]
  assign io_in_1_ready = grant_1 & io_out_ready; // @[Arbiter.scala 134:14]
  assign io_out_valid = _T_2 | io_in_1_valid; // @[Arbiter.scala 135:16]
  assign io_out_bits_setIdx = io_in_0_valid ? io_in_0_bits_setIdx : io_in_1_bits_setIdx; // @[Arbiter.scala 124:15 Arbiter.scala 128:19]
endmodule
module SRAMTemplateWithArbiter_5(
  input         clock,
  input         reset,
  output        io_r0_req_ready,
  input         io_r0_req_valid,
  input  [11:0] io_r0_req_bits_setIdx,
  output [63:0] io_r0_resp_data_0_data,
  output [63:0] io_r0_resp_data_1_data,
  output [63:0] io_r0_resp_data_2_data,
  output [63:0] io_r0_resp_data_3_data,
  output        io_r1_req_ready,
  input         io_r1_req_valid,
  input  [11:0] io_r1_req_bits_setIdx,
  output [63:0] io_r1_resp_data_0_data,
  output [63:0] io_r1_resp_data_1_data,
  output [63:0] io_r1_resp_data_2_data,
  output [63:0] io_r1_resp_data_3_data,
  input         io_wreq_valid,
  input  [11:0] io_wreq_bits_setIdx,
  input  [63:0] io_wreq_bits_data_data,
  input  [3:0]  io_wreq_bits_waymask
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [63:0] _RAND_1;
  reg [63:0] _RAND_2;
  reg [63:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [63:0] _RAND_8;
  reg [63:0] _RAND_9;
`endif // RANDOMIZE_REG_INIT
  wire  ram_clock; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rreq_ready; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_rreq_valid; // @[SRAMTemplate.scala 121:19]
  wire [11:0] ram_io_rreq_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_rresp_data_0_data; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_rresp_data_1_data; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_rresp_data_2_data; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_rresp_data_3_data; // @[SRAMTemplate.scala 121:19]
  wire  ram_io_wreq_valid; // @[SRAMTemplate.scala 121:19]
  wire [11:0] ram_io_wreq_bits_setIdx; // @[SRAMTemplate.scala 121:19]
  wire [63:0] ram_io_wreq_bits_data_data; // @[SRAMTemplate.scala 121:19]
  wire [3:0] ram_io_wreq_bits_waymask; // @[SRAMTemplate.scala 121:19]
  wire  readArb_io_in_0_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_0_valid; // @[SRAMTemplate.scala 124:23]
  wire [11:0] readArb_io_in_0_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_1_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_in_1_valid; // @[SRAMTemplate.scala 124:23]
  wire [11:0] readArb_io_in_1_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_ready; // @[SRAMTemplate.scala 124:23]
  wire  readArb_io_out_valid; // @[SRAMTemplate.scala 124:23]
  wire [11:0] readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 124:23]
  reg  _T_1; // @[SRAMTemplate.scala 130:58]
  reg [63:0] _T_3_0_data; // @[Reg.scala 27:20]
  reg [63:0] _T_3_1_data; // @[Reg.scala 27:20]
  reg [63:0] _T_3_2_data; // @[Reg.scala 27:20]
  reg [63:0] _T_3_3_data; // @[Reg.scala 27:20]
  reg  _T_6; // @[SRAMTemplate.scala 130:58]
  reg [63:0] _T_8_0_data; // @[Reg.scala 27:20]
  reg [63:0] _T_8_1_data; // @[Reg.scala 27:20]
  reg [63:0] _T_8_2_data; // @[Reg.scala 27:20]
  reg [63:0] _T_8_3_data; // @[Reg.scala 27:20]
  SRAMTemplate_6 ram ( // @[SRAMTemplate.scala 121:19]
    .clock(ram_clock),
    .io_rreq_ready(ram_io_rreq_ready),
    .io_rreq_valid(ram_io_rreq_valid),
    .io_rreq_bits_setIdx(ram_io_rreq_bits_setIdx),
    .io_rresp_data_0_data(ram_io_rresp_data_0_data),
    .io_rresp_data_1_data(ram_io_rresp_data_1_data),
    .io_rresp_data_2_data(ram_io_rresp_data_2_data),
    .io_rresp_data_3_data(ram_io_rresp_data_3_data),
    .io_wreq_valid(ram_io_wreq_valid),
    .io_wreq_bits_setIdx(ram_io_wreq_bits_setIdx),
    .io_wreq_bits_data_data(ram_io_wreq_bits_data_data),
    .io_wreq_bits_waymask(ram_io_wreq_bits_waymask)
  );
  Arbiter_13 readArb ( // @[SRAMTemplate.scala 124:23]
    .io_in_0_ready(readArb_io_in_0_ready),
    .io_in_0_valid(readArb_io_in_0_valid),
    .io_in_0_bits_setIdx(readArb_io_in_0_bits_setIdx),
    .io_in_1_ready(readArb_io_in_1_ready),
    .io_in_1_valid(readArb_io_in_1_valid),
    .io_in_1_bits_setIdx(readArb_io_in_1_bits_setIdx),
    .io_out_ready(readArb_io_out_ready),
    .io_out_valid(readArb_io_out_valid),
    .io_out_bits_setIdx(readArb_io_out_bits_setIdx)
  );
  assign io_r0_req_ready = readArb_io_in_0_ready; // @[SRAMTemplate.scala 125:17]
  assign io_r0_resp_data_0_data = _T_1 ? ram_io_rresp_data_0_data : _T_3_0_data; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_1_data = _T_1 ? ram_io_rresp_data_1_data : _T_3_1_data; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_2_data = _T_1 ? ram_io_rresp_data_2_data : _T_3_2_data; // @[SRAMTemplate.scala 130:17]
  assign io_r0_resp_data_3_data = _T_1 ? ram_io_rresp_data_3_data : _T_3_3_data; // @[SRAMTemplate.scala 130:17]
  assign io_r1_req_ready = readArb_io_in_1_ready; // @[SRAMTemplate.scala 125:17]
  assign io_r1_resp_data_0_data = _T_6 ? ram_io_rresp_data_0_data : _T_8_0_data; // @[SRAMTemplate.scala 130:17]
  assign io_r1_resp_data_1_data = _T_6 ? ram_io_rresp_data_1_data : _T_8_1_data; // @[SRAMTemplate.scala 130:17]
  assign io_r1_resp_data_2_data = _T_6 ? ram_io_rresp_data_2_data : _T_8_2_data; // @[SRAMTemplate.scala 130:17]
  assign io_r1_resp_data_3_data = _T_6 ? ram_io_rresp_data_3_data : _T_8_3_data; // @[SRAMTemplate.scala 130:17]
  assign ram_clock = clock;
  assign ram_io_rreq_valid = readArb_io_out_valid; // @[SRAMTemplate.scala 126:16]
  assign ram_io_rreq_bits_setIdx = readArb_io_out_bits_setIdx; // @[SRAMTemplate.scala 126:16]
  assign ram_io_wreq_valid = io_wreq_valid; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_setIdx = io_wreq_bits_setIdx; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_data_data = io_wreq_bits_data_data; // @[SRAMTemplate.scala 122:12]
  assign ram_io_wreq_bits_waymask = io_wreq_bits_waymask; // @[SRAMTemplate.scala 122:12]
  assign readArb_io_in_0_valid = io_r0_req_valid; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_0_bits_setIdx = io_r0_req_bits_setIdx; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_1_valid = io_r1_req_valid; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_in_1_bits_setIdx = io_r1_req_bits_setIdx; // @[SRAMTemplate.scala 125:17]
  assign readArb_io_out_ready = ram_io_rreq_ready; // @[SRAMTemplate.scala 126:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_1 = _RAND_0[0:0];
  _RAND_1 = {2{`RANDOM}};
  _T_3_0_data = _RAND_1[63:0];
  _RAND_2 = {2{`RANDOM}};
  _T_3_1_data = _RAND_2[63:0];
  _RAND_3 = {2{`RANDOM}};
  _T_3_2_data = _RAND_3[63:0];
  _RAND_4 = {2{`RANDOM}};
  _T_3_3_data = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  _T_6 = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  _T_8_0_data = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  _T_8_1_data = _RAND_7[63:0];
  _RAND_8 = {2{`RANDOM}};
  _T_8_2_data = _RAND_8[63:0];
  _RAND_9 = {2{`RANDOM}};
  _T_8_3_data = _RAND_9[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_1 <= io_r0_req_ready & io_r0_req_valid;
    if (reset) begin
      _T_3_0_data <= 64'h0;
    end else if (_T_1) begin
      _T_3_0_data <= ram_io_rresp_data_0_data;
    end
    if (reset) begin
      _T_3_1_data <= 64'h0;
    end else if (_T_1) begin
      _T_3_1_data <= ram_io_rresp_data_1_data;
    end
    if (reset) begin
      _T_3_2_data <= 64'h0;
    end else if (_T_1) begin
      _T_3_2_data <= ram_io_rresp_data_2_data;
    end
    if (reset) begin
      _T_3_3_data <= 64'h0;
    end else if (_T_1) begin
      _T_3_3_data <= ram_io_rresp_data_3_data;
    end
    _T_6 <= io_r1_req_ready & io_r1_req_valid;
    if (reset) begin
      _T_8_0_data <= 64'h0;
    end else if (_T_6) begin
      _T_8_0_data <= ram_io_rresp_data_0_data;
    end
    if (reset) begin
      _T_8_1_data <= 64'h0;
    end else if (_T_6) begin
      _T_8_1_data <= ram_io_rresp_data_1_data;
    end
    if (reset) begin
      _T_8_2_data <= 64'h0;
    end else if (_T_6) begin
      _T_8_2_data <= ram_io_rresp_data_2_data;
    end
    if (reset) begin
      _T_8_3_data <= 64'h0;
    end else if (_T_6) begin
      _T_8_3_data <= ram_io_rresp_data_3_data;
    end
  end
endmodule
module Cache_2(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_mem_req_ready,
  output        io_out_mem_req_valid,
  output [31:0] io_out_mem_req_bits_addr,
  output [3:0]  io_out_mem_req_bits_cmd,
  output [63:0] io_out_mem_req_bits_wdata,
  input         io_out_mem_resp_valid,
  input  [3:0]  io_out_mem_resp_bits_cmd,
  input  [63:0] io_out_mem_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [63:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [63:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [31:0] _RAND_21;
  reg [63:0] _RAND_22;
  reg [63:0] _RAND_23;
  reg [63:0] _RAND_24;
  reg [63:0] _RAND_25;
  reg [31:0] _RAND_26;
  reg [31:0] _RAND_27;
  reg [31:0] _RAND_28;
  reg [31:0] _RAND_29;
  reg [63:0] _RAND_30;
  reg [31:0] _RAND_31;
`endif // RANDOMIZE_REG_INIT
  wire  s1_io_in_ready; // @[Cache.scala 475:18]
  wire  s1_io_in_valid; // @[Cache.scala 475:18]
  wire [31:0] s1_io_in_bits_addr; // @[Cache.scala 475:18]
  wire [3:0] s1_io_in_bits_cmd; // @[Cache.scala 475:18]
  wire [7:0] s1_io_in_bits_wmask; // @[Cache.scala 475:18]
  wire [63:0] s1_io_in_bits_wdata; // @[Cache.scala 475:18]
  wire  s1_io_out_ready; // @[Cache.scala 475:18]
  wire  s1_io_out_valid; // @[Cache.scala 475:18]
  wire [31:0] s1_io_out_bits_req_addr; // @[Cache.scala 475:18]
  wire [3:0] s1_io_out_bits_req_cmd; // @[Cache.scala 475:18]
  wire [7:0] s1_io_out_bits_req_wmask; // @[Cache.scala 475:18]
  wire [63:0] s1_io_out_bits_req_wdata; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_req_ready; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_req_valid; // @[Cache.scala 475:18]
  wire [8:0] s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 475:18]
  wire [16:0] s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_0_dirty; // @[Cache.scala 475:18]
  wire [16:0] s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_1_dirty; // @[Cache.scala 475:18]
  wire [16:0] s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_2_dirty; // @[Cache.scala 475:18]
  wire [16:0] s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 475:18]
  wire  s1_io_metaReadBus_resp_data_3_dirty; // @[Cache.scala 475:18]
  wire  s1_io_dataReadBus_req_ready; // @[Cache.scala 475:18]
  wire  s1_io_dataReadBus_req_valid; // @[Cache.scala 475:18]
  wire [11:0] s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 475:18]
  wire [63:0] s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 475:18]
  wire [63:0] s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 475:18]
  wire [63:0] s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 475:18]
  wire [63:0] s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 475:18]
  wire  s2_clock; // @[Cache.scala 476:18]
  wire  s2_reset; // @[Cache.scala 476:18]
  wire  s2_io_in_ready; // @[Cache.scala 476:18]
  wire  s2_io_in_valid; // @[Cache.scala 476:18]
  wire [31:0] s2_io_in_bits_req_addr; // @[Cache.scala 476:18]
  wire [3:0] s2_io_in_bits_req_cmd; // @[Cache.scala 476:18]
  wire [7:0] s2_io_in_bits_req_wmask; // @[Cache.scala 476:18]
  wire [63:0] s2_io_in_bits_req_wdata; // @[Cache.scala 476:18]
  wire  s2_io_out_ready; // @[Cache.scala 476:18]
  wire  s2_io_out_valid; // @[Cache.scala 476:18]
  wire [31:0] s2_io_out_bits_req_addr; // @[Cache.scala 476:18]
  wire [3:0] s2_io_out_bits_req_cmd; // @[Cache.scala 476:18]
  wire [7:0] s2_io_out_bits_req_wmask; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_req_wdata; // @[Cache.scala 476:18]
  wire [16:0] s2_io_out_bits_metas_0_tag; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_0_valid; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_0_dirty; // @[Cache.scala 476:18]
  wire [16:0] s2_io_out_bits_metas_1_tag; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_1_valid; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_1_dirty; // @[Cache.scala 476:18]
  wire [16:0] s2_io_out_bits_metas_2_tag; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_2_valid; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_2_dirty; // @[Cache.scala 476:18]
  wire [16:0] s2_io_out_bits_metas_3_tag; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_3_valid; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_metas_3_dirty; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_datas_0_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_datas_1_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_datas_2_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_datas_3_data; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_hit; // @[Cache.scala 476:18]
  wire [3:0] s2_io_out_bits_waymask; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_mmio; // @[Cache.scala 476:18]
  wire  s2_io_out_bits_isForwardData; // @[Cache.scala 476:18]
  wire [63:0] s2_io_out_bits_forwardData_data_data; // @[Cache.scala 476:18]
  wire [3:0] s2_io_out_bits_forwardData_waymask; // @[Cache.scala 476:18]
  wire [16:0] s2_io_metaReadResp_0_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_0_valid; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_0_dirty; // @[Cache.scala 476:18]
  wire [16:0] s2_io_metaReadResp_1_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_1_valid; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_1_dirty; // @[Cache.scala 476:18]
  wire [16:0] s2_io_metaReadResp_2_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_2_valid; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_2_dirty; // @[Cache.scala 476:18]
  wire [16:0] s2_io_metaReadResp_3_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_3_valid; // @[Cache.scala 476:18]
  wire  s2_io_metaReadResp_3_dirty; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataReadResp_0_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataReadResp_1_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataReadResp_2_data; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataReadResp_3_data; // @[Cache.scala 476:18]
  wire  s2_io_metaWriteBus_req_valid; // @[Cache.scala 476:18]
  wire [8:0] s2_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 476:18]
  wire [16:0] s2_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 476:18]
  wire  s2_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 476:18]
  wire [3:0] s2_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 476:18]
  wire  s2_io_dataWriteBus_req_valid; // @[Cache.scala 476:18]
  wire [11:0] s2_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 476:18]
  wire [63:0] s2_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 476:18]
  wire [3:0] s2_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 476:18]
  wire  s3_clock; // @[Cache.scala 477:18]
  wire  s3_reset; // @[Cache.scala 477:18]
  wire  s3_io_in_ready; // @[Cache.scala 477:18]
  wire  s3_io_in_valid; // @[Cache.scala 477:18]
  wire [31:0] s3_io_in_bits_req_addr; // @[Cache.scala 477:18]
  wire [3:0] s3_io_in_bits_req_cmd; // @[Cache.scala 477:18]
  wire [7:0] s3_io_in_bits_req_wmask; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_req_wdata; // @[Cache.scala 477:18]
  wire [16:0] s3_io_in_bits_metas_0_tag; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_0_valid; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_0_dirty; // @[Cache.scala 477:18]
  wire [16:0] s3_io_in_bits_metas_1_tag; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_1_valid; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_1_dirty; // @[Cache.scala 477:18]
  wire [16:0] s3_io_in_bits_metas_2_tag; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_2_valid; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_2_dirty; // @[Cache.scala 477:18]
  wire [16:0] s3_io_in_bits_metas_3_tag; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_3_valid; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_metas_3_dirty; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_datas_0_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_datas_1_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_datas_2_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_datas_3_data; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_hit; // @[Cache.scala 477:18]
  wire [3:0] s3_io_in_bits_waymask; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_mmio; // @[Cache.scala 477:18]
  wire  s3_io_in_bits_isForwardData; // @[Cache.scala 477:18]
  wire [63:0] s3_io_in_bits_forwardData_data_data; // @[Cache.scala 477:18]
  wire [3:0] s3_io_in_bits_forwardData_waymask; // @[Cache.scala 477:18]
  wire  s3_io_out_valid; // @[Cache.scala 477:18]
  wire [3:0] s3_io_out_bits_cmd; // @[Cache.scala 477:18]
  wire [63:0] s3_io_out_bits_rdata; // @[Cache.scala 477:18]
  wire  s3_io_isFinish; // @[Cache.scala 477:18]
  wire  s3_io_dataReadBus_req_ready; // @[Cache.scala 477:18]
  wire  s3_io_dataReadBus_req_valid; // @[Cache.scala 477:18]
  wire [11:0] s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataReadBus_resp_data_0_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataReadBus_resp_data_1_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataReadBus_resp_data_2_data; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataReadBus_resp_data_3_data; // @[Cache.scala 477:18]
  wire  s3_io_dataWriteBus_req_valid; // @[Cache.scala 477:18]
  wire [11:0] s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 477:18]
  wire [63:0] s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 477:18]
  wire [3:0] s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 477:18]
  wire  s3_io_metaWriteBus_req_valid; // @[Cache.scala 477:18]
  wire [8:0] s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 477:18]
  wire [16:0] s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 477:18]
  wire  s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 477:18]
  wire [3:0] s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 477:18]
  wire  s3_io_mem_req_ready; // @[Cache.scala 477:18]
  wire  s3_io_mem_req_valid; // @[Cache.scala 477:18]
  wire [31:0] s3_io_mem_req_bits_addr; // @[Cache.scala 477:18]
  wire [3:0] s3_io_mem_req_bits_cmd; // @[Cache.scala 477:18]
  wire [63:0] s3_io_mem_req_bits_wdata; // @[Cache.scala 477:18]
  wire  s3_io_mem_resp_ready; // @[Cache.scala 477:18]
  wire  s3_io_mem_resp_valid; // @[Cache.scala 477:18]
  wire [3:0] s3_io_mem_resp_bits_cmd; // @[Cache.scala 477:18]
  wire [63:0] s3_io_mem_resp_bits_rdata; // @[Cache.scala 477:18]
  wire  s3_io_cohResp_valid; // @[Cache.scala 477:18]
  wire  s3_io_dataReadRespToL1; // @[Cache.scala 477:18]
  wire  metaArray_clock; // @[Cache.scala 478:25]
  wire  metaArray_reset; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_req_ready; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_req_valid; // @[Cache.scala 478:25]
  wire [8:0] metaArray_io_r0_req_bits_setIdx; // @[Cache.scala 478:25]
  wire [16:0] metaArray_io_r0_resp_data_0_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_resp_data_0_valid; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_resp_data_0_dirty; // @[Cache.scala 478:25]
  wire [16:0] metaArray_io_r0_resp_data_1_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_resp_data_1_valid; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_resp_data_1_dirty; // @[Cache.scala 478:25]
  wire [16:0] metaArray_io_r0_resp_data_2_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_resp_data_2_valid; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_resp_data_2_dirty; // @[Cache.scala 478:25]
  wire [16:0] metaArray_io_r0_resp_data_3_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_resp_data_3_valid; // @[Cache.scala 478:25]
  wire  metaArray_io_r0_resp_data_3_dirty; // @[Cache.scala 478:25]
  wire  metaArray_io_wreq_valid; // @[Cache.scala 478:25]
  wire [8:0] metaArray_io_wreq_bits_setIdx; // @[Cache.scala 478:25]
  wire [16:0] metaArray_io_wreq_bits_data_tag; // @[Cache.scala 478:25]
  wire  metaArray_io_wreq_bits_data_dirty; // @[Cache.scala 478:25]
  wire [3:0] metaArray_io_wreq_bits_waymask; // @[Cache.scala 478:25]
  wire  dataArray_clock; // @[Cache.scala 479:25]
  wire  dataArray_reset; // @[Cache.scala 479:25]
  wire  dataArray_io_r0_req_ready; // @[Cache.scala 479:25]
  wire  dataArray_io_r0_req_valid; // @[Cache.scala 479:25]
  wire [11:0] dataArray_io_r0_req_bits_setIdx; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r0_resp_data_0_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r0_resp_data_1_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r0_resp_data_2_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r0_resp_data_3_data; // @[Cache.scala 479:25]
  wire  dataArray_io_r1_req_ready; // @[Cache.scala 479:25]
  wire  dataArray_io_r1_req_valid; // @[Cache.scala 479:25]
  wire [11:0] dataArray_io_r1_req_bits_setIdx; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r1_resp_data_0_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r1_resp_data_1_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r1_resp_data_2_data; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_r1_resp_data_3_data; // @[Cache.scala 479:25]
  wire  dataArray_io_wreq_valid; // @[Cache.scala 479:25]
  wire [11:0] dataArray_io_wreq_bits_setIdx; // @[Cache.scala 479:25]
  wire [63:0] dataArray_io_wreq_bits_data_data; // @[Cache.scala 479:25]
  wire [3:0] dataArray_io_wreq_bits_waymask; // @[Cache.scala 479:25]
  wire  arb_io_in_0_ready; // @[Cache.scala 488:19]
  wire  arb_io_in_0_valid; // @[Cache.scala 488:19]
  wire [31:0] arb_io_in_0_bits_addr; // @[Cache.scala 488:19]
  wire [2:0] arb_io_in_0_bits_size; // @[Cache.scala 488:19]
  wire [3:0] arb_io_in_0_bits_cmd; // @[Cache.scala 488:19]
  wire [7:0] arb_io_in_0_bits_wmask; // @[Cache.scala 488:19]
  wire [63:0] arb_io_in_0_bits_wdata; // @[Cache.scala 488:19]
  wire  arb_io_in_1_ready; // @[Cache.scala 488:19]
  wire  arb_io_in_1_valid; // @[Cache.scala 488:19]
  wire [31:0] arb_io_in_1_bits_addr; // @[Cache.scala 488:19]
  wire [2:0] arb_io_in_1_bits_size; // @[Cache.scala 488:19]
  wire [3:0] arb_io_in_1_bits_cmd; // @[Cache.scala 488:19]
  wire [7:0] arb_io_in_1_bits_wmask; // @[Cache.scala 488:19]
  wire [63:0] arb_io_in_1_bits_wdata; // @[Cache.scala 488:19]
  wire  arb_io_out_ready; // @[Cache.scala 488:19]
  wire  arb_io_out_valid; // @[Cache.scala 488:19]
  wire [31:0] arb_io_out_bits_addr; // @[Cache.scala 488:19]
  wire [2:0] arb_io_out_bits_size; // @[Cache.scala 488:19]
  wire [3:0] arb_io_out_bits_cmd; // @[Cache.scala 488:19]
  wire [7:0] arb_io_out_bits_wmask; // @[Cache.scala 488:19]
  wire [63:0] arb_io_out_bits_wdata; // @[Cache.scala 488:19]
  wire  _T = s2_io_out_ready & s2_io_out_valid; // @[Decoupled.scala 40:37]
  reg  _T_2; // @[Pipeline.scala 24:24]
  wire  _GEN_0 = _T ? 1'h0 : _T_2; // @[Pipeline.scala 25:25]
  wire  _T_3 = s1_io_out_valid & s2_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_1 = _T_3 | _GEN_0; // @[Pipeline.scala 26:38]
  reg [31:0] _T_5_req_addr; // @[Reg.scala 15:16]
  reg [3:0] _T_5_req_cmd; // @[Reg.scala 15:16]
  reg [7:0] _T_5_req_wmask; // @[Reg.scala 15:16]
  reg [63:0] _T_5_req_wdata; // @[Reg.scala 15:16]
  reg  _T_7; // @[Pipeline.scala 24:24]
  wire  _GEN_8 = s3_io_isFinish ? 1'h0 : _T_7; // @[Pipeline.scala 25:25]
  wire  _T_8 = s2_io_out_valid & s3_io_in_ready; // @[Pipeline.scala 26:22]
  wire  _GEN_9 = _T_8 | _GEN_8; // @[Pipeline.scala 26:38]
  reg [31:0] _T_10_req_addr; // @[Reg.scala 15:16]
  reg [3:0] _T_10_req_cmd; // @[Reg.scala 15:16]
  reg [7:0] _T_10_req_wmask; // @[Reg.scala 15:16]
  reg [63:0] _T_10_req_wdata; // @[Reg.scala 15:16]
  reg [16:0] _T_10_metas_0_tag; // @[Reg.scala 15:16]
  reg  _T_10_metas_0_valid; // @[Reg.scala 15:16]
  reg  _T_10_metas_0_dirty; // @[Reg.scala 15:16]
  reg [16:0] _T_10_metas_1_tag; // @[Reg.scala 15:16]
  reg  _T_10_metas_1_valid; // @[Reg.scala 15:16]
  reg  _T_10_metas_1_dirty; // @[Reg.scala 15:16]
  reg [16:0] _T_10_metas_2_tag; // @[Reg.scala 15:16]
  reg  _T_10_metas_2_valid; // @[Reg.scala 15:16]
  reg  _T_10_metas_2_dirty; // @[Reg.scala 15:16]
  reg [16:0] _T_10_metas_3_tag; // @[Reg.scala 15:16]
  reg  _T_10_metas_3_valid; // @[Reg.scala 15:16]
  reg  _T_10_metas_3_dirty; // @[Reg.scala 15:16]
  reg [63:0] _T_10_datas_0_data; // @[Reg.scala 15:16]
  reg [63:0] _T_10_datas_1_data; // @[Reg.scala 15:16]
  reg [63:0] _T_10_datas_2_data; // @[Reg.scala 15:16]
  reg [63:0] _T_10_datas_3_data; // @[Reg.scala 15:16]
  reg  _T_10_hit; // @[Reg.scala 15:16]
  reg [3:0] _T_10_waymask; // @[Reg.scala 15:16]
  reg  _T_10_mmio; // @[Reg.scala 15:16]
  reg  _T_10_isForwardData; // @[Reg.scala 15:16]
  reg [63:0] _T_10_forwardData_data_data; // @[Reg.scala 15:16]
  reg [3:0] _T_10_forwardData_waymask; // @[Reg.scala 15:16]
  wire  _T_15 = s3_io_out_bits_cmd == 4'h4; // @[SimpleBus.scala 95:26]
  wire  _T_16 = s3_io_out_valid & _T_15; // @[Cache.scala 505:43]
  wire  _T_17 = s3_io_out_valid | s3_io_dataReadRespToL1; // @[Cache.scala 505:100]
  CacheStage1_2 s1 ( // @[Cache.scala 475:18]
    .io_in_ready(s1_io_in_ready),
    .io_in_valid(s1_io_in_valid),
    .io_in_bits_addr(s1_io_in_bits_addr),
    .io_in_bits_cmd(s1_io_in_bits_cmd),
    .io_in_bits_wmask(s1_io_in_bits_wmask),
    .io_in_bits_wdata(s1_io_in_bits_wdata),
    .io_out_ready(s1_io_out_ready),
    .io_out_valid(s1_io_out_valid),
    .io_out_bits_req_addr(s1_io_out_bits_req_addr),
    .io_out_bits_req_cmd(s1_io_out_bits_req_cmd),
    .io_out_bits_req_wmask(s1_io_out_bits_req_wmask),
    .io_out_bits_req_wdata(s1_io_out_bits_req_wdata),
    .io_metaReadBus_req_ready(s1_io_metaReadBus_req_ready),
    .io_metaReadBus_req_valid(s1_io_metaReadBus_req_valid),
    .io_metaReadBus_req_bits_setIdx(s1_io_metaReadBus_req_bits_setIdx),
    .io_metaReadBus_resp_data_0_tag(s1_io_metaReadBus_resp_data_0_tag),
    .io_metaReadBus_resp_data_0_valid(s1_io_metaReadBus_resp_data_0_valid),
    .io_metaReadBus_resp_data_0_dirty(s1_io_metaReadBus_resp_data_0_dirty),
    .io_metaReadBus_resp_data_1_tag(s1_io_metaReadBus_resp_data_1_tag),
    .io_metaReadBus_resp_data_1_valid(s1_io_metaReadBus_resp_data_1_valid),
    .io_metaReadBus_resp_data_1_dirty(s1_io_metaReadBus_resp_data_1_dirty),
    .io_metaReadBus_resp_data_2_tag(s1_io_metaReadBus_resp_data_2_tag),
    .io_metaReadBus_resp_data_2_valid(s1_io_metaReadBus_resp_data_2_valid),
    .io_metaReadBus_resp_data_2_dirty(s1_io_metaReadBus_resp_data_2_dirty),
    .io_metaReadBus_resp_data_3_tag(s1_io_metaReadBus_resp_data_3_tag),
    .io_metaReadBus_resp_data_3_valid(s1_io_metaReadBus_resp_data_3_valid),
    .io_metaReadBus_resp_data_3_dirty(s1_io_metaReadBus_resp_data_3_dirty),
    .io_dataReadBus_req_ready(s1_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s1_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s1_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s1_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s1_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s1_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s1_io_dataReadBus_resp_data_3_data)
  );
  CacheStage2_2 s2 ( // @[Cache.scala 476:18]
    .clock(s2_clock),
    .reset(s2_reset),
    .io_in_ready(s2_io_in_ready),
    .io_in_valid(s2_io_in_valid),
    .io_in_bits_req_addr(s2_io_in_bits_req_addr),
    .io_in_bits_req_cmd(s2_io_in_bits_req_cmd),
    .io_in_bits_req_wmask(s2_io_in_bits_req_wmask),
    .io_in_bits_req_wdata(s2_io_in_bits_req_wdata),
    .io_out_ready(s2_io_out_ready),
    .io_out_valid(s2_io_out_valid),
    .io_out_bits_req_addr(s2_io_out_bits_req_addr),
    .io_out_bits_req_cmd(s2_io_out_bits_req_cmd),
    .io_out_bits_req_wmask(s2_io_out_bits_req_wmask),
    .io_out_bits_req_wdata(s2_io_out_bits_req_wdata),
    .io_out_bits_metas_0_tag(s2_io_out_bits_metas_0_tag),
    .io_out_bits_metas_0_valid(s2_io_out_bits_metas_0_valid),
    .io_out_bits_metas_0_dirty(s2_io_out_bits_metas_0_dirty),
    .io_out_bits_metas_1_tag(s2_io_out_bits_metas_1_tag),
    .io_out_bits_metas_1_valid(s2_io_out_bits_metas_1_valid),
    .io_out_bits_metas_1_dirty(s2_io_out_bits_metas_1_dirty),
    .io_out_bits_metas_2_tag(s2_io_out_bits_metas_2_tag),
    .io_out_bits_metas_2_valid(s2_io_out_bits_metas_2_valid),
    .io_out_bits_metas_2_dirty(s2_io_out_bits_metas_2_dirty),
    .io_out_bits_metas_3_tag(s2_io_out_bits_metas_3_tag),
    .io_out_bits_metas_3_valid(s2_io_out_bits_metas_3_valid),
    .io_out_bits_metas_3_dirty(s2_io_out_bits_metas_3_dirty),
    .io_out_bits_datas_0_data(s2_io_out_bits_datas_0_data),
    .io_out_bits_datas_1_data(s2_io_out_bits_datas_1_data),
    .io_out_bits_datas_2_data(s2_io_out_bits_datas_2_data),
    .io_out_bits_datas_3_data(s2_io_out_bits_datas_3_data),
    .io_out_bits_hit(s2_io_out_bits_hit),
    .io_out_bits_waymask(s2_io_out_bits_waymask),
    .io_out_bits_mmio(s2_io_out_bits_mmio),
    .io_out_bits_isForwardData(s2_io_out_bits_isForwardData),
    .io_out_bits_forwardData_data_data(s2_io_out_bits_forwardData_data_data),
    .io_out_bits_forwardData_waymask(s2_io_out_bits_forwardData_waymask),
    .io_metaReadResp_0_tag(s2_io_metaReadResp_0_tag),
    .io_metaReadResp_0_valid(s2_io_metaReadResp_0_valid),
    .io_metaReadResp_0_dirty(s2_io_metaReadResp_0_dirty),
    .io_metaReadResp_1_tag(s2_io_metaReadResp_1_tag),
    .io_metaReadResp_1_valid(s2_io_metaReadResp_1_valid),
    .io_metaReadResp_1_dirty(s2_io_metaReadResp_1_dirty),
    .io_metaReadResp_2_tag(s2_io_metaReadResp_2_tag),
    .io_metaReadResp_2_valid(s2_io_metaReadResp_2_valid),
    .io_metaReadResp_2_dirty(s2_io_metaReadResp_2_dirty),
    .io_metaReadResp_3_tag(s2_io_metaReadResp_3_tag),
    .io_metaReadResp_3_valid(s2_io_metaReadResp_3_valid),
    .io_metaReadResp_3_dirty(s2_io_metaReadResp_3_dirty),
    .io_dataReadResp_0_data(s2_io_dataReadResp_0_data),
    .io_dataReadResp_1_data(s2_io_dataReadResp_1_data),
    .io_dataReadResp_2_data(s2_io_dataReadResp_2_data),
    .io_dataReadResp_3_data(s2_io_dataReadResp_3_data),
    .io_metaWriteBus_req_valid(s2_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s2_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s2_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_dirty(s2_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s2_io_metaWriteBus_req_bits_waymask),
    .io_dataWriteBus_req_valid(s2_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s2_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s2_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s2_io_dataWriteBus_req_bits_waymask)
  );
  CacheStage3_2 s3 ( // @[Cache.scala 477:18]
    .clock(s3_clock),
    .reset(s3_reset),
    .io_in_ready(s3_io_in_ready),
    .io_in_valid(s3_io_in_valid),
    .io_in_bits_req_addr(s3_io_in_bits_req_addr),
    .io_in_bits_req_cmd(s3_io_in_bits_req_cmd),
    .io_in_bits_req_wmask(s3_io_in_bits_req_wmask),
    .io_in_bits_req_wdata(s3_io_in_bits_req_wdata),
    .io_in_bits_metas_0_tag(s3_io_in_bits_metas_0_tag),
    .io_in_bits_metas_0_valid(s3_io_in_bits_metas_0_valid),
    .io_in_bits_metas_0_dirty(s3_io_in_bits_metas_0_dirty),
    .io_in_bits_metas_1_tag(s3_io_in_bits_metas_1_tag),
    .io_in_bits_metas_1_valid(s3_io_in_bits_metas_1_valid),
    .io_in_bits_metas_1_dirty(s3_io_in_bits_metas_1_dirty),
    .io_in_bits_metas_2_tag(s3_io_in_bits_metas_2_tag),
    .io_in_bits_metas_2_valid(s3_io_in_bits_metas_2_valid),
    .io_in_bits_metas_2_dirty(s3_io_in_bits_metas_2_dirty),
    .io_in_bits_metas_3_tag(s3_io_in_bits_metas_3_tag),
    .io_in_bits_metas_3_valid(s3_io_in_bits_metas_3_valid),
    .io_in_bits_metas_3_dirty(s3_io_in_bits_metas_3_dirty),
    .io_in_bits_datas_0_data(s3_io_in_bits_datas_0_data),
    .io_in_bits_datas_1_data(s3_io_in_bits_datas_1_data),
    .io_in_bits_datas_2_data(s3_io_in_bits_datas_2_data),
    .io_in_bits_datas_3_data(s3_io_in_bits_datas_3_data),
    .io_in_bits_hit(s3_io_in_bits_hit),
    .io_in_bits_waymask(s3_io_in_bits_waymask),
    .io_in_bits_mmio(s3_io_in_bits_mmio),
    .io_in_bits_isForwardData(s3_io_in_bits_isForwardData),
    .io_in_bits_forwardData_data_data(s3_io_in_bits_forwardData_data_data),
    .io_in_bits_forwardData_waymask(s3_io_in_bits_forwardData_waymask),
    .io_out_valid(s3_io_out_valid),
    .io_out_bits_cmd(s3_io_out_bits_cmd),
    .io_out_bits_rdata(s3_io_out_bits_rdata),
    .io_isFinish(s3_io_isFinish),
    .io_dataReadBus_req_ready(s3_io_dataReadBus_req_ready),
    .io_dataReadBus_req_valid(s3_io_dataReadBus_req_valid),
    .io_dataReadBus_req_bits_setIdx(s3_io_dataReadBus_req_bits_setIdx),
    .io_dataReadBus_resp_data_0_data(s3_io_dataReadBus_resp_data_0_data),
    .io_dataReadBus_resp_data_1_data(s3_io_dataReadBus_resp_data_1_data),
    .io_dataReadBus_resp_data_2_data(s3_io_dataReadBus_resp_data_2_data),
    .io_dataReadBus_resp_data_3_data(s3_io_dataReadBus_resp_data_3_data),
    .io_dataWriteBus_req_valid(s3_io_dataWriteBus_req_valid),
    .io_dataWriteBus_req_bits_setIdx(s3_io_dataWriteBus_req_bits_setIdx),
    .io_dataWriteBus_req_bits_data_data(s3_io_dataWriteBus_req_bits_data_data),
    .io_dataWriteBus_req_bits_waymask(s3_io_dataWriteBus_req_bits_waymask),
    .io_metaWriteBus_req_valid(s3_io_metaWriteBus_req_valid),
    .io_metaWriteBus_req_bits_setIdx(s3_io_metaWriteBus_req_bits_setIdx),
    .io_metaWriteBus_req_bits_data_tag(s3_io_metaWriteBus_req_bits_data_tag),
    .io_metaWriteBus_req_bits_data_dirty(s3_io_metaWriteBus_req_bits_data_dirty),
    .io_metaWriteBus_req_bits_waymask(s3_io_metaWriteBus_req_bits_waymask),
    .io_mem_req_ready(s3_io_mem_req_ready),
    .io_mem_req_valid(s3_io_mem_req_valid),
    .io_mem_req_bits_addr(s3_io_mem_req_bits_addr),
    .io_mem_req_bits_cmd(s3_io_mem_req_bits_cmd),
    .io_mem_req_bits_wdata(s3_io_mem_req_bits_wdata),
    .io_mem_resp_ready(s3_io_mem_resp_ready),
    .io_mem_resp_valid(s3_io_mem_resp_valid),
    .io_mem_resp_bits_cmd(s3_io_mem_resp_bits_cmd),
    .io_mem_resp_bits_rdata(s3_io_mem_resp_bits_rdata),
    .io_cohResp_valid(s3_io_cohResp_valid),
    .io_dataReadRespToL1(s3_io_dataReadRespToL1)
  );
  SRAMTemplateWithArbiter_4 metaArray ( // @[Cache.scala 478:25]
    .clock(metaArray_clock),
    .reset(metaArray_reset),
    .io_r0_req_ready(metaArray_io_r0_req_ready),
    .io_r0_req_valid(metaArray_io_r0_req_valid),
    .io_r0_req_bits_setIdx(metaArray_io_r0_req_bits_setIdx),
    .io_r0_resp_data_0_tag(metaArray_io_r0_resp_data_0_tag),
    .io_r0_resp_data_0_valid(metaArray_io_r0_resp_data_0_valid),
    .io_r0_resp_data_0_dirty(metaArray_io_r0_resp_data_0_dirty),
    .io_r0_resp_data_1_tag(metaArray_io_r0_resp_data_1_tag),
    .io_r0_resp_data_1_valid(metaArray_io_r0_resp_data_1_valid),
    .io_r0_resp_data_1_dirty(metaArray_io_r0_resp_data_1_dirty),
    .io_r0_resp_data_2_tag(metaArray_io_r0_resp_data_2_tag),
    .io_r0_resp_data_2_valid(metaArray_io_r0_resp_data_2_valid),
    .io_r0_resp_data_2_dirty(metaArray_io_r0_resp_data_2_dirty),
    .io_r0_resp_data_3_tag(metaArray_io_r0_resp_data_3_tag),
    .io_r0_resp_data_3_valid(metaArray_io_r0_resp_data_3_valid),
    .io_r0_resp_data_3_dirty(metaArray_io_r0_resp_data_3_dirty),
    .io_wreq_valid(metaArray_io_wreq_valid),
    .io_wreq_bits_setIdx(metaArray_io_wreq_bits_setIdx),
    .io_wreq_bits_data_tag(metaArray_io_wreq_bits_data_tag),
    .io_wreq_bits_data_dirty(metaArray_io_wreq_bits_data_dirty),
    .io_wreq_bits_waymask(metaArray_io_wreq_bits_waymask)
  );
  SRAMTemplateWithArbiter_5 dataArray ( // @[Cache.scala 479:25]
    .clock(dataArray_clock),
    .reset(dataArray_reset),
    .io_r0_req_ready(dataArray_io_r0_req_ready),
    .io_r0_req_valid(dataArray_io_r0_req_valid),
    .io_r0_req_bits_setIdx(dataArray_io_r0_req_bits_setIdx),
    .io_r0_resp_data_0_data(dataArray_io_r0_resp_data_0_data),
    .io_r0_resp_data_1_data(dataArray_io_r0_resp_data_1_data),
    .io_r0_resp_data_2_data(dataArray_io_r0_resp_data_2_data),
    .io_r0_resp_data_3_data(dataArray_io_r0_resp_data_3_data),
    .io_r1_req_ready(dataArray_io_r1_req_ready),
    .io_r1_req_valid(dataArray_io_r1_req_valid),
    .io_r1_req_bits_setIdx(dataArray_io_r1_req_bits_setIdx),
    .io_r1_resp_data_0_data(dataArray_io_r1_resp_data_0_data),
    .io_r1_resp_data_1_data(dataArray_io_r1_resp_data_1_data),
    .io_r1_resp_data_2_data(dataArray_io_r1_resp_data_2_data),
    .io_r1_resp_data_3_data(dataArray_io_r1_resp_data_3_data),
    .io_wreq_valid(dataArray_io_wreq_valid),
    .io_wreq_bits_setIdx(dataArray_io_wreq_bits_setIdx),
    .io_wreq_bits_data_data(dataArray_io_wreq_bits_data_data),
    .io_wreq_bits_waymask(dataArray_io_wreq_bits_waymask)
  );
  Arbiter_9 arb ( // @[Cache.scala 488:19]
    .io_in_0_ready(arb_io_in_0_ready),
    .io_in_0_valid(arb_io_in_0_valid),
    .io_in_0_bits_addr(arb_io_in_0_bits_addr),
    .io_in_0_bits_size(arb_io_in_0_bits_size),
    .io_in_0_bits_cmd(arb_io_in_0_bits_cmd),
    .io_in_0_bits_wmask(arb_io_in_0_bits_wmask),
    .io_in_0_bits_wdata(arb_io_in_0_bits_wdata),
    .io_in_1_ready(arb_io_in_1_ready),
    .io_in_1_valid(arb_io_in_1_valid),
    .io_in_1_bits_addr(arb_io_in_1_bits_addr),
    .io_in_1_bits_size(arb_io_in_1_bits_size),
    .io_in_1_bits_cmd(arb_io_in_1_bits_cmd),
    .io_in_1_bits_wmask(arb_io_in_1_bits_wmask),
    .io_in_1_bits_wdata(arb_io_in_1_bits_wdata),
    .io_out_ready(arb_io_out_ready),
    .io_out_valid(arb_io_out_valid),
    .io_out_bits_addr(arb_io_out_bits_addr),
    .io_out_bits_size(arb_io_out_bits_size),
    .io_out_bits_cmd(arb_io_out_bits_cmd),
    .io_out_bits_wmask(arb_io_out_bits_wmask),
    .io_out_bits_wdata(arb_io_out_bits_wdata)
  );
  assign io_in_req_ready = arb_io_in_1_ready; // @[Cache.scala 489:28]
  assign io_in_resp_valid = _T_16 ? 1'h0 : _T_17; // @[Cache.scala 499:14 Cache.scala 505:20]
  assign io_in_resp_bits_cmd = s3_io_out_bits_cmd; // @[Cache.scala 499:14]
  assign io_in_resp_bits_rdata = s3_io_out_bits_rdata; // @[Cache.scala 499:14]
  assign io_out_mem_req_valid = s3_io_mem_req_valid; // @[Cache.scala 501:14]
  assign io_out_mem_req_bits_addr = s3_io_mem_req_bits_addr; // @[Cache.scala 501:14]
  assign io_out_mem_req_bits_cmd = s3_io_mem_req_bits_cmd; // @[Cache.scala 501:14]
  assign io_out_mem_req_bits_wdata = s3_io_mem_req_bits_wdata; // @[Cache.scala 501:14]
  assign s1_io_in_valid = arb_io_out_valid; // @[Cache.scala 491:12]
  assign s1_io_in_bits_addr = arb_io_out_bits_addr; // @[Cache.scala 491:12]
  assign s1_io_in_bits_cmd = arb_io_out_bits_cmd; // @[Cache.scala 491:12]
  assign s1_io_in_bits_wmask = arb_io_out_bits_wmask; // @[Cache.scala 491:12]
  assign s1_io_in_bits_wdata = arb_io_out_bits_wdata; // @[Cache.scala 491:12]
  assign s1_io_out_ready = s2_io_in_ready; // @[Pipeline.scala 29:16]
  assign s1_io_metaReadBus_req_ready = metaArray_io_r0_req_ready; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_0_tag = metaArray_io_r0_resp_data_0_tag; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_0_valid = metaArray_io_r0_resp_data_0_valid; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_0_dirty = metaArray_io_r0_resp_data_0_dirty; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_1_tag = metaArray_io_r0_resp_data_1_tag; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_1_valid = metaArray_io_r0_resp_data_1_valid; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_1_dirty = metaArray_io_r0_resp_data_1_dirty; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_2_tag = metaArray_io_r0_resp_data_2_tag; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_2_valid = metaArray_io_r0_resp_data_2_valid; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_2_dirty = metaArray_io_r0_resp_data_2_dirty; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_3_tag = metaArray_io_r0_resp_data_3_tag; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_3_valid = metaArray_io_r0_resp_data_3_valid; // @[Cache.scala 523:21]
  assign s1_io_metaReadBus_resp_data_3_dirty = metaArray_io_r0_resp_data_3_dirty; // @[Cache.scala 523:21]
  assign s1_io_dataReadBus_req_ready = dataArray_io_r0_req_ready; // @[Cache.scala 524:21]
  assign s1_io_dataReadBus_resp_data_0_data = dataArray_io_r0_resp_data_0_data; // @[Cache.scala 524:21]
  assign s1_io_dataReadBus_resp_data_1_data = dataArray_io_r0_resp_data_1_data; // @[Cache.scala 524:21]
  assign s1_io_dataReadBus_resp_data_2_data = dataArray_io_r0_resp_data_2_data; // @[Cache.scala 524:21]
  assign s1_io_dataReadBus_resp_data_3_data = dataArray_io_r0_resp_data_3_data; // @[Cache.scala 524:21]
  assign s2_clock = clock;
  assign s2_reset = reset;
  assign s2_io_in_valid = _T_2; // @[Pipeline.scala 31:17]
  assign s2_io_in_bits_req_addr = _T_5_req_addr; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_cmd = _T_5_req_cmd; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_wmask = _T_5_req_wmask; // @[Pipeline.scala 30:16]
  assign s2_io_in_bits_req_wdata = _T_5_req_wdata; // @[Pipeline.scala 30:16]
  assign s2_io_out_ready = s3_io_in_ready; // @[Pipeline.scala 29:16]
  assign s2_io_metaReadResp_0_tag = s1_io_metaReadBus_resp_data_0_tag; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_0_valid = s1_io_metaReadBus_resp_data_0_valid; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_0_dirty = s1_io_metaReadBus_resp_data_0_dirty; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_1_tag = s1_io_metaReadBus_resp_data_1_tag; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_1_valid = s1_io_metaReadBus_resp_data_1_valid; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_1_dirty = s1_io_metaReadBus_resp_data_1_dirty; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_2_tag = s1_io_metaReadBus_resp_data_2_tag; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_2_valid = s1_io_metaReadBus_resp_data_2_valid; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_2_dirty = s1_io_metaReadBus_resp_data_2_dirty; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_3_tag = s1_io_metaReadBus_resp_data_3_tag; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_3_valid = s1_io_metaReadBus_resp_data_3_valid; // @[Cache.scala 530:22]
  assign s2_io_metaReadResp_3_dirty = s1_io_metaReadBus_resp_data_3_dirty; // @[Cache.scala 530:22]
  assign s2_io_dataReadResp_0_data = s1_io_dataReadBus_resp_data_0_data; // @[Cache.scala 531:22]
  assign s2_io_dataReadResp_1_data = s1_io_dataReadBus_resp_data_1_data; // @[Cache.scala 531:22]
  assign s2_io_dataReadResp_2_data = s1_io_dataReadBus_resp_data_2_data; // @[Cache.scala 531:22]
  assign s2_io_dataReadResp_3_data = s1_io_dataReadBus_resp_data_3_data; // @[Cache.scala 531:22]
  assign s2_io_metaWriteBus_req_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 533:22]
  assign s2_io_metaWriteBus_req_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 533:22]
  assign s2_io_metaWriteBus_req_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 533:22]
  assign s2_io_metaWriteBus_req_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 533:22]
  assign s2_io_metaWriteBus_req_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 533:22]
  assign s2_io_dataWriteBus_req_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 532:22]
  assign s2_io_dataWriteBus_req_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 532:22]
  assign s2_io_dataWriteBus_req_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 532:22]
  assign s2_io_dataWriteBus_req_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 532:22]
  assign s3_clock = clock;
  assign s3_reset = reset;
  assign s3_io_in_valid = _T_7; // @[Pipeline.scala 31:17]
  assign s3_io_in_bits_req_addr = _T_10_req_addr; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_cmd = _T_10_req_cmd; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_wmask = _T_10_req_wmask; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_req_wdata = _T_10_req_wdata; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_tag = _T_10_metas_0_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_valid = _T_10_metas_0_valid; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_0_dirty = _T_10_metas_0_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_tag = _T_10_metas_1_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_valid = _T_10_metas_1_valid; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_1_dirty = _T_10_metas_1_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_tag = _T_10_metas_2_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_valid = _T_10_metas_2_valid; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_2_dirty = _T_10_metas_2_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_tag = _T_10_metas_3_tag; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_valid = _T_10_metas_3_valid; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_metas_3_dirty = _T_10_metas_3_dirty; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_0_data = _T_10_datas_0_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_1_data = _T_10_datas_1_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_2_data = _T_10_datas_2_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_datas_3_data = _T_10_datas_3_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_hit = _T_10_hit; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_waymask = _T_10_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_mmio = _T_10_mmio; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_isForwardData = _T_10_isForwardData; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_data_data = _T_10_forwardData_data_data; // @[Pipeline.scala 30:16]
  assign s3_io_in_bits_forwardData_waymask = _T_10_forwardData_waymask; // @[Pipeline.scala 30:16]
  assign s3_io_dataReadBus_req_ready = dataArray_io_r1_req_ready; // @[Cache.scala 525:21]
  assign s3_io_dataReadBus_resp_data_0_data = dataArray_io_r1_resp_data_0_data; // @[Cache.scala 525:21]
  assign s3_io_dataReadBus_resp_data_1_data = dataArray_io_r1_resp_data_1_data; // @[Cache.scala 525:21]
  assign s3_io_dataReadBus_resp_data_2_data = dataArray_io_r1_resp_data_2_data; // @[Cache.scala 525:21]
  assign s3_io_dataReadBus_resp_data_3_data = dataArray_io_r1_resp_data_3_data; // @[Cache.scala 525:21]
  assign s3_io_mem_req_ready = io_out_mem_req_ready; // @[Cache.scala 501:14]
  assign s3_io_mem_resp_valid = io_out_mem_resp_valid; // @[Cache.scala 501:14]
  assign s3_io_mem_resp_bits_cmd = io_out_mem_resp_bits_cmd; // @[Cache.scala 501:14]
  assign s3_io_mem_resp_bits_rdata = io_out_mem_resp_bits_rdata; // @[Cache.scala 501:14]
  assign metaArray_clock = clock;
  assign metaArray_reset = reset;
  assign metaArray_io_r0_req_valid = s1_io_metaReadBus_req_valid; // @[Cache.scala 523:21]
  assign metaArray_io_r0_req_bits_setIdx = s1_io_metaReadBus_req_bits_setIdx; // @[Cache.scala 523:21]
  assign metaArray_io_wreq_valid = s3_io_metaWriteBus_req_valid; // @[Cache.scala 527:18]
  assign metaArray_io_wreq_bits_setIdx = s3_io_metaWriteBus_req_bits_setIdx; // @[Cache.scala 527:18]
  assign metaArray_io_wreq_bits_data_tag = s3_io_metaWriteBus_req_bits_data_tag; // @[Cache.scala 527:18]
  assign metaArray_io_wreq_bits_data_dirty = s3_io_metaWriteBus_req_bits_data_dirty; // @[Cache.scala 527:18]
  assign metaArray_io_wreq_bits_waymask = s3_io_metaWriteBus_req_bits_waymask; // @[Cache.scala 527:18]
  assign dataArray_clock = clock;
  assign dataArray_reset = reset;
  assign dataArray_io_r0_req_valid = s1_io_dataReadBus_req_valid; // @[Cache.scala 524:21]
  assign dataArray_io_r0_req_bits_setIdx = s1_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 524:21]
  assign dataArray_io_r1_req_valid = s3_io_dataReadBus_req_valid; // @[Cache.scala 525:21]
  assign dataArray_io_r1_req_bits_setIdx = s3_io_dataReadBus_req_bits_setIdx; // @[Cache.scala 525:21]
  assign dataArray_io_wreq_valid = s3_io_dataWriteBus_req_valid; // @[Cache.scala 528:18]
  assign dataArray_io_wreq_bits_setIdx = s3_io_dataWriteBus_req_bits_setIdx; // @[Cache.scala 528:18]
  assign dataArray_io_wreq_bits_data_data = s3_io_dataWriteBus_req_bits_data_data; // @[Cache.scala 528:18]
  assign dataArray_io_wreq_bits_waymask = s3_io_dataWriteBus_req_bits_waymask; // @[Cache.scala 528:18]
  assign arb_io_in_0_valid = 1'h0; // @[Cache.scala 513:24]
  assign arb_io_in_0_bits_addr = 32'h0; // @[Cache.scala 512:23]
  assign arb_io_in_0_bits_size = 3'h0; // @[Cache.scala 512:23]
  assign arb_io_in_0_bits_cmd = 4'h0; // @[Cache.scala 512:23]
  assign arb_io_in_0_bits_wmask = 8'h0; // @[Cache.scala 512:23]
  assign arb_io_in_0_bits_wdata = 64'h0; // @[Cache.scala 512:23]
  assign arb_io_in_1_valid = io_in_req_valid; // @[Cache.scala 489:28]
  assign arb_io_in_1_bits_addr = io_in_req_bits_addr; // @[Cache.scala 489:28]
  assign arb_io_in_1_bits_size = io_in_req_bits_size; // @[Cache.scala 489:28]
  assign arb_io_in_1_bits_cmd = io_in_req_bits_cmd; // @[Cache.scala 489:28]
  assign arb_io_in_1_bits_wmask = io_in_req_bits_wmask; // @[Cache.scala 489:28]
  assign arb_io_in_1_bits_wdata = io_in_req_bits_wdata; // @[Cache.scala 489:28]
  assign arb_io_out_ready = s1_io_in_ready; // @[Cache.scala 491:12]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  _T_5_req_addr = _RAND_1[31:0];
  _RAND_2 = {1{`RANDOM}};
  _T_5_req_cmd = _RAND_2[3:0];
  _RAND_3 = {1{`RANDOM}};
  _T_5_req_wmask = _RAND_3[7:0];
  _RAND_4 = {2{`RANDOM}};
  _T_5_req_wdata = _RAND_4[63:0];
  _RAND_5 = {1{`RANDOM}};
  _T_7 = _RAND_5[0:0];
  _RAND_6 = {1{`RANDOM}};
  _T_10_req_addr = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  _T_10_req_cmd = _RAND_7[3:0];
  _RAND_8 = {1{`RANDOM}};
  _T_10_req_wmask = _RAND_8[7:0];
  _RAND_9 = {2{`RANDOM}};
  _T_10_req_wdata = _RAND_9[63:0];
  _RAND_10 = {1{`RANDOM}};
  _T_10_metas_0_tag = _RAND_10[16:0];
  _RAND_11 = {1{`RANDOM}};
  _T_10_metas_0_valid = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _T_10_metas_0_dirty = _RAND_12[0:0];
  _RAND_13 = {1{`RANDOM}};
  _T_10_metas_1_tag = _RAND_13[16:0];
  _RAND_14 = {1{`RANDOM}};
  _T_10_metas_1_valid = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  _T_10_metas_1_dirty = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  _T_10_metas_2_tag = _RAND_16[16:0];
  _RAND_17 = {1{`RANDOM}};
  _T_10_metas_2_valid = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _T_10_metas_2_dirty = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  _T_10_metas_3_tag = _RAND_19[16:0];
  _RAND_20 = {1{`RANDOM}};
  _T_10_metas_3_valid = _RAND_20[0:0];
  _RAND_21 = {1{`RANDOM}};
  _T_10_metas_3_dirty = _RAND_21[0:0];
  _RAND_22 = {2{`RANDOM}};
  _T_10_datas_0_data = _RAND_22[63:0];
  _RAND_23 = {2{`RANDOM}};
  _T_10_datas_1_data = _RAND_23[63:0];
  _RAND_24 = {2{`RANDOM}};
  _T_10_datas_2_data = _RAND_24[63:0];
  _RAND_25 = {2{`RANDOM}};
  _T_10_datas_3_data = _RAND_25[63:0];
  _RAND_26 = {1{`RANDOM}};
  _T_10_hit = _RAND_26[0:0];
  _RAND_27 = {1{`RANDOM}};
  _T_10_waymask = _RAND_27[3:0];
  _RAND_28 = {1{`RANDOM}};
  _T_10_mmio = _RAND_28[0:0];
  _RAND_29 = {1{`RANDOM}};
  _T_10_isForwardData = _RAND_29[0:0];
  _RAND_30 = {2{`RANDOM}};
  _T_10_forwardData_data_data = _RAND_30[63:0];
  _RAND_31 = {1{`RANDOM}};
  _T_10_forwardData_waymask = _RAND_31[3:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_2 <= 1'h0;
    end else begin
      _T_2 <= _GEN_1;
    end
    if (_T_3) begin
      _T_5_req_addr <= s1_io_out_bits_req_addr;
    end
    if (_T_3) begin
      _T_5_req_cmd <= s1_io_out_bits_req_cmd;
    end
    if (_T_3) begin
      _T_5_req_wmask <= s1_io_out_bits_req_wmask;
    end
    if (_T_3) begin
      _T_5_req_wdata <= s1_io_out_bits_req_wdata;
    end
    if (reset) begin
      _T_7 <= 1'h0;
    end else begin
      _T_7 <= _GEN_9;
    end
    if (_T_8) begin
      _T_10_req_addr <= s2_io_out_bits_req_addr;
    end
    if (_T_8) begin
      _T_10_req_cmd <= s2_io_out_bits_req_cmd;
    end
    if (_T_8) begin
      _T_10_req_wmask <= s2_io_out_bits_req_wmask;
    end
    if (_T_8) begin
      _T_10_req_wdata <= s2_io_out_bits_req_wdata;
    end
    if (_T_8) begin
      _T_10_metas_0_tag <= s2_io_out_bits_metas_0_tag;
    end
    if (_T_8) begin
      _T_10_metas_0_valid <= s2_io_out_bits_metas_0_valid;
    end
    if (_T_8) begin
      _T_10_metas_0_dirty <= s2_io_out_bits_metas_0_dirty;
    end
    if (_T_8) begin
      _T_10_metas_1_tag <= s2_io_out_bits_metas_1_tag;
    end
    if (_T_8) begin
      _T_10_metas_1_valid <= s2_io_out_bits_metas_1_valid;
    end
    if (_T_8) begin
      _T_10_metas_1_dirty <= s2_io_out_bits_metas_1_dirty;
    end
    if (_T_8) begin
      _T_10_metas_2_tag <= s2_io_out_bits_metas_2_tag;
    end
    if (_T_8) begin
      _T_10_metas_2_valid <= s2_io_out_bits_metas_2_valid;
    end
    if (_T_8) begin
      _T_10_metas_2_dirty <= s2_io_out_bits_metas_2_dirty;
    end
    if (_T_8) begin
      _T_10_metas_3_tag <= s2_io_out_bits_metas_3_tag;
    end
    if (_T_8) begin
      _T_10_metas_3_valid <= s2_io_out_bits_metas_3_valid;
    end
    if (_T_8) begin
      _T_10_metas_3_dirty <= s2_io_out_bits_metas_3_dirty;
    end
    if (_T_8) begin
      _T_10_datas_0_data <= s2_io_out_bits_datas_0_data;
    end
    if (_T_8) begin
      _T_10_datas_1_data <= s2_io_out_bits_datas_1_data;
    end
    if (_T_8) begin
      _T_10_datas_2_data <= s2_io_out_bits_datas_2_data;
    end
    if (_T_8) begin
      _T_10_datas_3_data <= s2_io_out_bits_datas_3_data;
    end
    if (_T_8) begin
      _T_10_hit <= s2_io_out_bits_hit;
    end
    if (_T_8) begin
      _T_10_waymask <= s2_io_out_bits_waymask;
    end
    if (_T_8) begin
      _T_10_mmio <= s2_io_out_bits_mmio;
    end
    if (_T_8) begin
      _T_10_isForwardData <= s2_io_out_bits_isForwardData;
    end
    if (_T_8) begin
      _T_10_forwardData_data_data <= s2_io_out_bits_forwardData_data_data;
    end
    if (_T_8) begin
      _T_10_forwardData_waymask <= s2_io_out_bits_forwardData_waymask;
    end
  end
endmodule
module SimpleBusAddressMapper(
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [3:0]  io_in_req_bits_cmd,
  input  [63:0] io_in_req_bits_wdata,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_req_ready,
  output        io_out_req_valid,
  output [31:0] io_out_req_bits_addr,
  output [3:0]  io_out_req_bits_cmd,
  output [63:0] io_out_req_bits_wdata,
  input         io_out_resp_valid,
  input  [3:0]  io_out_resp_bits_cmd,
  input  [63:0] io_out_resp_bits_rdata
);
  assign io_in_req_ready = io_out_req_ready; // @[AddressMapper.scala 31:10]
  assign io_in_resp_valid = io_out_resp_valid; // @[AddressMapper.scala 31:10]
  assign io_in_resp_bits_cmd = io_out_resp_bits_cmd; // @[AddressMapper.scala 31:10]
  assign io_in_resp_bits_rdata = io_out_resp_bits_rdata; // @[AddressMapper.scala 31:10]
  assign io_out_req_valid = io_in_req_valid; // @[AddressMapper.scala 31:10]
  assign io_out_req_bits_addr = {4'h1,io_in_req_bits_addr[27:0]}; // @[AddressMapper.scala 31:10 AddressMapper.scala 34:26]
  assign io_out_req_bits_cmd = io_in_req_bits_cmd; // @[AddressMapper.scala 31:10]
  assign io_out_req_bits_wdata = io_in_req_bits_wdata; // @[AddressMapper.scala 31:10]
endmodule
module SimpleBus2AXI4Converter(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [3:0]  io_in_req_bits_cmd,
  input  [63:0] io_in_req_bits_wdata,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_awready,
  output        io_out_awvalid,
  output [31:0] io_out_awaddr,
  output [2:0]  io_out_awprot,
  output        io_out_awid,
  output        io_out_awuser,
  output [7:0]  io_out_awlen,
  output [2:0]  io_out_awsize,
  output [1:0]  io_out_awburst,
  output        io_out_awlock,
  output [3:0]  io_out_awcache,
  output [3:0]  io_out_awqos,
  input         io_out_wready,
  output        io_out_wvalid,
  output [63:0] io_out_wdata,
  output        io_out_wlast,
  input         io_out_bvalid,
  input         io_out_arready,
  output        io_out_arvalid,
  output [31:0] io_out_araddr,
  output [2:0]  io_out_arprot,
  output        io_out_arid,
  output        io_out_aruser,
  output [7:0]  io_out_arlen,
  output [2:0]  io_out_arsize,
  output [1:0]  io_out_arburst,
  output        io_out_arlock,
  output [3:0]  io_out_arcache,
  output [3:0]  io_out_arqos,
  input         io_out_rvalid,
  input  [63:0] io_out_rdata,
  input         io_out_rlast
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] _T_8 = io_in_req_bits_cmd[1] ? 3'h7 : 3'h0; // @[ToAXI4.scala 169:30]
  wire  _T_9 = io_in_req_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_10 = io_in_req_bits_cmd == 4'h1; // @[SimpleBus.scala 77:29]
  wire [2:0] _T_12 = io_out_rlast ? 3'h6 : 3'h0; // @[ToAXI4.scala 184:28]
  wire  _T_13 = io_out_awready & io_out_awvalid; // @[Decoupled.scala 40:37]
  reg  awAck; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_13 | awAck; // @[StopWatch.scala 30:20]
  wire  _T_17 = io_out_wready & io_out_wvalid; // @[Decoupled.scala 40:37]
  wire  _T_18 = _T_13 & _T_17; // @[ToAXI4.scala 189:27]
  wire  _T_19 = _T_18 & io_out_wlast; // @[ToAXI4.scala 189:43]
  reg  wAck; // @[StopWatch.scala 24:20]
  wire  _T_20 = awAck & wAck; // @[ToAXI4.scala 189:63]
  wire  wSend = _T_19 | _T_20; // @[ToAXI4.scala 189:53]
  wire  _T_15 = _T_17 & io_out_wlast; // @[ToAXI4.scala 188:41]
  wire  _GEN_2 = _T_15 | wAck; // @[StopWatch.scala 30:20]
  wire  _T_23 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 40:37]
  reg  wen; // @[Reg.scala 15:16]
  wire  _T_25 = ~io_in_req_bits_cmd[0]; // @[SimpleBus.scala 73:18]
  wire  _T_27 = ~io_in_req_bits_cmd[3]; // @[SimpleBus.scala 73:29]
  wire  _T_28 = _T_25 & _T_27; // @[SimpleBus.scala 73:26]
  wire  _T_31 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[SimpleBus.scala 103:29]
  wire  _T_32 = ~awAck; // @[ToAXI4.scala 193:36]
  wire  _T_36 = ~wAck; // @[ToAXI4.scala 194:36]
  wire  _T_40 = _T_36 & io_out_wready; // @[ToAXI4.scala 195:55]
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _T_40 : io_out_arready; // @[ToAXI4.scala 195:18]
  assign io_in_resp_valid = wen ? io_out_bvalid : io_out_rvalid; // @[ToAXI4.scala 199:19]
  assign io_in_resp_bits_cmd = {{1'd0}, _T_12}; // @[ToAXI4.scala 184:22]
  assign io_in_resp_bits_rdata = io_out_rdata; // @[ToAXI4.scala 183:23]
  assign io_out_awvalid = _T_31 & _T_32; // @[ToAXI4.scala 193:16]
  assign io_out_awaddr = io_out_araddr; // @[ToAXI4.scala 182:6]
  assign io_out_awprot = io_out_arprot; // @[ToAXI4.scala 182:6]
  assign io_out_awid = io_out_arid; // @[ToAXI4.scala 182:6]
  assign io_out_awuser = io_out_aruser; // @[ToAXI4.scala 182:6]
  assign io_out_awlen = io_out_arlen; // @[ToAXI4.scala 182:6]
  assign io_out_awsize = io_out_arsize; // @[ToAXI4.scala 182:6]
  assign io_out_awburst = io_out_arburst; // @[ToAXI4.scala 182:6]
  assign io_out_awlock = io_out_arlock; // @[ToAXI4.scala 182:6]
  assign io_out_awcache = io_out_arcache; // @[ToAXI4.scala 182:6]
  assign io_out_awqos = io_out_arqos; // @[ToAXI4.scala 182:6]
  assign io_out_wvalid = _T_31 & _T_36; // @[ToAXI4.scala 194:16]
  assign io_out_wdata = io_in_req_bits_wdata; // @[ToAXI4.scala 160:10]
  assign io_out_wlast = _T_9 | _T_10; // @[ToAXI4.scala 177:24]
  assign io_out_arvalid = io_in_req_valid & _T_28; // @[ToAXI4.scala 192:16]
  assign io_out_araddr = io_in_req_bits_addr; // @[ToAXI4.scala 158:12]
  assign io_out_arprot = 3'h1; // @[ToAXI4.scala 159:12]
  assign io_out_arid = 1'h0; // @[ToAXI4.scala 168:24]
  assign io_out_aruser = 1'h0; // @[ToAXI4.scala 176:24]
  assign io_out_arlen = {{5'd0}, _T_8}; // @[ToAXI4.scala 169:24]
  assign io_out_arsize = 3'h3; // @[ToAXI4.scala 170:24]
  assign io_out_arburst = 2'h2; // @[ToAXI4.scala 171:24]
  assign io_out_arlock = 1'h0; // @[ToAXI4.scala 173:24]
  assign io_out_arcache = 4'h0; // @[ToAXI4.scala 174:24]
  assign io_out_arqos = 4'h0; // @[ToAXI4.scala 175:24]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  awAck = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wen = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      awAck <= 1'h0;
    end else if (wSend) begin
      awAck <= 1'h0;
    end else begin
      awAck <= _GEN_0;
    end
    if (reset) begin
      wAck <= 1'h0;
    end else if (wSend) begin
      wAck <= 1'h0;
    end else begin
      wAck <= _GEN_2;
    end
    if (_T_23) begin
      wen <= io_in_req_bits_cmd[0];
    end
  end
endmodule
module SimpleBusCrossbar1toN(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_0_req_ready,
  output        io_out_0_req_valid,
  output [31:0] io_out_0_req_bits_addr,
  output [2:0]  io_out_0_req_bits_size,
  output [3:0]  io_out_0_req_bits_cmd,
  output [7:0]  io_out_0_req_bits_wmask,
  output [63:0] io_out_0_req_bits_wdata,
  output        io_out_0_resp_ready,
  input         io_out_0_resp_valid,
  input  [3:0]  io_out_0_resp_bits_cmd,
  input  [63:0] io_out_0_resp_bits_rdata,
  input         io_out_1_req_ready,
  output        io_out_1_req_valid,
  output [31:0] io_out_1_req_bits_addr,
  output [3:0]  io_out_1_req_bits_cmd,
  output [7:0]  io_out_1_req_bits_wmask,
  output [63:0] io_out_1_req_bits_wdata,
  output        io_out_1_resp_ready,
  input         io_out_1_resp_valid,
  input  [63:0] io_out_1_resp_bits_rdata,
  input         io_out_2_req_ready,
  output        io_out_2_req_valid,
  output [31:0] io_out_2_req_bits_addr,
  output [3:0]  io_out_2_req_bits_cmd,
  output [7:0]  io_out_2_req_bits_wmask,
  output [63:0] io_out_2_req_bits_wdata,
  output        io_out_2_resp_ready,
  input         io_out_2_resp_valid,
  input  [63:0] io_out_2_resp_bits_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  reg [1:0] state; // @[Crossbar.scala 31:22]
  wire  outSelVec_0 = io_in_req_bits_addr >= 32'he0000000; // @[Crossbar.scala 36:20]
  wire  _T_3 = io_in_req_bits_addr >= 32'h38000000; // @[Crossbar.scala 36:20]
  wire  _T_4 = io_in_req_bits_addr < 32'h38010000; // @[Crossbar.scala 36:42]
  wire  outSelVec_1 = _T_3 & _T_4; // @[Crossbar.scala 36:34]
  wire  _T_6 = io_in_req_bits_addr >= 32'h3c000000; // @[Crossbar.scala 36:20]
  wire  _T_7 = io_in_req_bits_addr < 32'h40000000; // @[Crossbar.scala 36:42]
  wire  outSelVec_2 = _T_6 & _T_7; // @[Crossbar.scala 36:34]
  wire [1:0] _T_9 = outSelVec_1 ? 2'h1 : 2'h2; // @[Mux.scala 47:69]
  wire [1:0] outSelIdx = outSelVec_0 ? 2'h0 : _T_9; // @[Mux.scala 47:69]
  wire  _GEN_11 = 2'h1 == outSelIdx ? io_out_1_req_ready : io_out_0_req_ready; // @[Decoupled.scala 40:37]
  wire  _GEN_12 = 2'h1 == outSelIdx ? io_out_1_req_valid : io_out_0_req_valid; // @[Decoupled.scala 40:37]
  wire  _GEN_22 = 2'h2 == outSelIdx ? io_out_2_req_ready : _GEN_11; // @[Decoupled.scala 40:37]
  wire  _GEN_23 = 2'h2 == outSelIdx ? io_out_2_req_valid : _GEN_12; // @[Decoupled.scala 40:37]
  wire  _T_10 = _GEN_22 & _GEN_23; // @[Decoupled.scala 40:37]
  wire  _T_11 = state == 2'h0; // @[Crossbar.scala 39:72]
  wire  _T_12 = _T_10 & _T_11; // @[Crossbar.scala 39:62]
  reg [1:0] outSelIdxResp; // @[Reg.scala 15:16]
  wire [2:0] _T_14 = {outSelVec_2,outSelVec_1,outSelVec_0}; // @[Crossbar.scala 41:54]
  wire  _T_15 = |_T_14; // @[Crossbar.scala 41:61]
  wire  _T_16 = ~_T_15; // @[Crossbar.scala 41:43]
  wire  reqInvalidAddr = io_in_req_valid & _T_16; // @[Crossbar.scala 41:40]
  wire  _T_24 = &_T_14; // @[Crossbar.scala 43:91]
  wire  _T_25 = io_in_req_valid & _T_24; // @[Crossbar.scala 43:71]
  wire  _T_38 = ~_T_25; // @[Crossbar.scala 49:10]
  wire  _T_40 = _T_38 | reset; // @[Crossbar.scala 49:9]
  wire  _T_41 = ~_T_40; // @[Crossbar.scala 49:9]
  wire  _T_43 = io_in_req_valid & _T_11; // @[Crossbar.scala 54:42]
  wire  _T_51 = 2'h0 == state; // @[Conditional.scala 37:30]
  wire  _T_53 = 2'h1 == state; // @[Conditional.scala 37:30]
  wire  _GEN_54 = 2'h1 == outSelIdxResp ? io_out_1_resp_ready : io_out_0_resp_ready; // @[Decoupled.scala 40:37]
  wire  _GEN_55 = 2'h1 == outSelIdxResp ? io_out_1_resp_valid : io_out_0_resp_valid; // @[Decoupled.scala 40:37]
  wire [3:0] _GEN_56 = 2'h1 == outSelIdxResp ? 4'h6 : io_out_0_resp_bits_cmd; // @[Decoupled.scala 40:37]
  wire [63:0] _GEN_57 = 2'h1 == outSelIdxResp ? io_out_1_resp_bits_rdata : io_out_0_resp_bits_rdata; // @[Decoupled.scala 40:37]
  wire  _GEN_65 = 2'h2 == outSelIdxResp ? io_out_2_resp_ready : _GEN_54; // @[Decoupled.scala 40:37]
  wire  _GEN_66 = 2'h2 == outSelIdxResp ? io_out_2_resp_valid : _GEN_55; // @[Decoupled.scala 40:37]
  wire  _T_54 = _GEN_65 & _GEN_66; // @[Decoupled.scala 40:37]
  wire  _T_55 = 2'h2 == state; // @[Conditional.scala 37:30]
  wire  _T_58 = state == 2'h2; // @[Crossbar.scala 67:55]
  wire  _GEN_77 = 2'h0 == outSelIdxResp; // @[Crossbar.scala 70:25]
  wire  _GEN_78 = 2'h1 == outSelIdxResp; // @[Crossbar.scala 70:25]
  wire  _GEN_79 = 2'h2 == outSelIdxResp; // @[Crossbar.scala 70:25]
  assign io_in_req_ready = _GEN_22 | reqInvalidAddr; // @[Crossbar.scala 71:19]
  assign io_in_resp_valid = _T_54 | _T_58; // @[Crossbar.scala 67:20]
  assign io_in_resp_bits_cmd = 2'h2 == outSelIdxResp ? 4'h6 : _GEN_56; // @[Crossbar.scala 68:19]
  assign io_in_resp_bits_rdata = 2'h2 == outSelIdxResp ? io_out_2_resp_bits_rdata : _GEN_57; // @[Crossbar.scala 68:19]
  assign io_out_0_req_valid = outSelVec_0 & _T_43; // @[Crossbar.scala 54:17]
  assign io_out_0_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 53:16]
  assign io_out_0_req_bits_size = io_in_req_bits_size; // @[Crossbar.scala 53:16]
  assign io_out_0_req_bits_cmd = io_in_req_bits_cmd; // @[Crossbar.scala 53:16]
  assign io_out_0_req_bits_wmask = io_in_req_bits_wmask; // @[Crossbar.scala 53:16]
  assign io_out_0_req_bits_wdata = io_in_req_bits_wdata; // @[Crossbar.scala 53:16]
  assign io_out_0_resp_ready = _GEN_77 | outSelVec_0; // @[Crossbar.scala 55:18 Crossbar.scala 70:25]
  assign io_out_1_req_valid = outSelVec_1 & _T_43; // @[Crossbar.scala 54:17]
  assign io_out_1_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 53:16]
  assign io_out_1_req_bits_cmd = io_in_req_bits_cmd; // @[Crossbar.scala 53:16]
  assign io_out_1_req_bits_wmask = io_in_req_bits_wmask; // @[Crossbar.scala 53:16]
  assign io_out_1_req_bits_wdata = io_in_req_bits_wdata; // @[Crossbar.scala 53:16]
  assign io_out_1_resp_ready = _GEN_78 | outSelVec_1; // @[Crossbar.scala 55:18 Crossbar.scala 70:25]
  assign io_out_2_req_valid = outSelVec_2 & _T_43; // @[Crossbar.scala 54:17]
  assign io_out_2_req_bits_addr = io_in_req_bits_addr; // @[Crossbar.scala 53:16]
  assign io_out_2_req_bits_cmd = io_in_req_bits_cmd; // @[Crossbar.scala 53:16]
  assign io_out_2_req_bits_wmask = io_in_req_bits_wmask; // @[Crossbar.scala 53:16]
  assign io_out_2_req_bits_wdata = io_in_req_bits_wdata; // @[Crossbar.scala 53:16]
  assign io_out_2_resp_ready = _GEN_79 | outSelVec_2; // @[Crossbar.scala 55:18 Crossbar.scala 70:25]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  _RAND_1 = {1{`RANDOM}};
  outSelIdxResp = _RAND_1[1:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else if (_T_51) begin
      if (reqInvalidAddr) begin
        state <= 2'h2;
      end else if (_T_10) begin
        state <= 2'h1;
      end
    end else if (_T_53) begin
      if (_T_54) begin
        state <= 2'h0;
      end
    end else if (_T_55) begin
      if (io_in_resp_valid) begin
        state <= 2'h0;
      end
    end
    if (_T_12) begin
      if (outSelVec_0) begin
        outSelIdxResp <= 2'h0;
      end else if (outSelVec_1) begin
        outSelIdxResp <= 2'h1;
      end else begin
        outSelIdxResp <= 2'h2;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_41) begin
          $fwrite(32'h80000002,"Assertion failed: address decode error, bad addr = 0x%x\n\n    at Crossbar.scala:49 assert(!(io.in.req.valid && outSelVec.asUInt.andR), \"address decode error, bad addr = 0x%%x\\n\", addr)\n",io_in_req_bits_addr); // @[Crossbar.scala 49:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_41) begin
          $fatal; // @[Crossbar.scala 49:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module SimpleBus2AXI4Converter_1(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [2:0]  io_in_req_bits_size,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [3:0]  io_in_resp_bits_cmd,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_awready,
  output        io_out_awvalid,
  output [31:0] io_out_awaddr,
  output [2:0]  io_out_awprot,
  output        io_out_awid,
  output        io_out_awuser,
  output [7:0]  io_out_awlen,
  output [2:0]  io_out_awsize,
  output [1:0]  io_out_awburst,
  output        io_out_awlock,
  output [3:0]  io_out_awcache,
  output [3:0]  io_out_awqos,
  input         io_out_wready,
  output        io_out_wvalid,
  output [63:0] io_out_wdata,
  output [7:0]  io_out_wstrb,
  output        io_out_wlast,
  output        io_out_bready,
  input         io_out_bvalid,
  input         io_out_arready,
  output        io_out_arvalid,
  output [31:0] io_out_araddr,
  output [2:0]  io_out_arprot,
  output        io_out_arid,
  output        io_out_aruser,
  output [7:0]  io_out_arlen,
  output [2:0]  io_out_arsize,
  output [1:0]  io_out_arburst,
  output        io_out_arlock,
  output [3:0]  io_out_arcache,
  output [3:0]  io_out_arqos,
  output        io_out_rready,
  input         io_out_rvalid,
  input  [63:0] io_out_rdata,
  input         io_out_rlast
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire [2:0] _T_8 = io_in_req_bits_cmd[1] ? 3'h7 : 3'h0; // @[ToAXI4.scala 169:30]
  wire  _T_9 = io_in_req_bits_cmd == 4'h7; // @[SimpleBus.scala 78:27]
  wire  _T_10 = io_in_req_bits_cmd == 4'h1; // @[SimpleBus.scala 77:29]
  wire [2:0] _T_12 = io_out_rlast ? 3'h6 : 3'h0; // @[ToAXI4.scala 184:28]
  wire  _T_13 = io_out_awready & io_out_awvalid; // @[Decoupled.scala 40:37]
  reg  awAck; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_13 | awAck; // @[StopWatch.scala 30:20]
  wire  _T_17 = io_out_wready & io_out_wvalid; // @[Decoupled.scala 40:37]
  wire  _T_18 = _T_13 & _T_17; // @[ToAXI4.scala 189:27]
  wire  _T_19 = _T_18 & io_out_wlast; // @[ToAXI4.scala 189:43]
  reg  wAck; // @[StopWatch.scala 24:20]
  wire  _T_20 = awAck & wAck; // @[ToAXI4.scala 189:63]
  wire  wSend = _T_19 | _T_20; // @[ToAXI4.scala 189:53]
  wire  _T_15 = _T_17 & io_out_wlast; // @[ToAXI4.scala 188:41]
  wire  _GEN_2 = _T_15 | wAck; // @[StopWatch.scala 30:20]
  wire  _T_23 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 40:37]
  reg  wen; // @[Reg.scala 15:16]
  wire  _T_25 = ~io_in_req_bits_cmd[0]; // @[SimpleBus.scala 73:18]
  wire  _T_27 = ~io_in_req_bits_cmd[3]; // @[SimpleBus.scala 73:29]
  wire  _T_28 = _T_25 & _T_27; // @[SimpleBus.scala 73:26]
  wire  _T_31 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[SimpleBus.scala 103:29]
  wire  _T_32 = ~awAck; // @[ToAXI4.scala 193:36]
  wire  _T_36 = ~wAck; // @[ToAXI4.scala 194:36]
  wire  _T_40 = _T_36 & io_out_wready; // @[ToAXI4.scala 195:55]
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _T_40 : io_out_arready; // @[ToAXI4.scala 195:18]
  assign io_in_resp_valid = wen ? io_out_bvalid : io_out_rvalid; // @[ToAXI4.scala 199:19]
  assign io_in_resp_bits_cmd = {{1'd0}, _T_12}; // @[ToAXI4.scala 184:22]
  assign io_in_resp_bits_rdata = io_out_rdata; // @[ToAXI4.scala 183:23]
  assign io_out_awvalid = _T_31 & _T_32; // @[ToAXI4.scala 193:16]
  assign io_out_awaddr = io_out_araddr; // @[ToAXI4.scala 182:6]
  assign io_out_awprot = io_out_arprot; // @[ToAXI4.scala 182:6]
  assign io_out_awid = io_out_arid; // @[ToAXI4.scala 182:6]
  assign io_out_awuser = io_out_aruser; // @[ToAXI4.scala 182:6]
  assign io_out_awlen = io_out_arlen; // @[ToAXI4.scala 182:6]
  assign io_out_awsize = io_out_arsize; // @[ToAXI4.scala 182:6]
  assign io_out_awburst = io_out_arburst; // @[ToAXI4.scala 182:6]
  assign io_out_awlock = io_out_arlock; // @[ToAXI4.scala 182:6]
  assign io_out_awcache = io_out_arcache; // @[ToAXI4.scala 182:6]
  assign io_out_awqos = io_out_arqos; // @[ToAXI4.scala 182:6]
  assign io_out_wvalid = _T_31 & _T_36; // @[ToAXI4.scala 194:16]
  assign io_out_wdata = io_in_req_bits_wdata; // @[ToAXI4.scala 160:10]
  assign io_out_wstrb = io_in_req_bits_wmask; // @[ToAXI4.scala 161:10]
  assign io_out_wlast = _T_9 | _T_10; // @[ToAXI4.scala 177:24]
  assign io_out_bready = io_in_resp_ready; // @[ToAXI4.scala 198:16]
  assign io_out_arvalid = io_in_req_valid & _T_28; // @[ToAXI4.scala 192:16]
  assign io_out_araddr = io_in_req_bits_addr; // @[ToAXI4.scala 158:12]
  assign io_out_arprot = 3'h1; // @[ToAXI4.scala 159:12]
  assign io_out_arid = 1'h0; // @[ToAXI4.scala 168:24]
  assign io_out_aruser = 1'h0; // @[ToAXI4.scala 176:24]
  assign io_out_arlen = {{5'd0}, _T_8}; // @[ToAXI4.scala 169:24]
  assign io_out_arsize = io_in_req_bits_size; // @[ToAXI4.scala 170:24]
  assign io_out_arburst = 2'h1; // @[ToAXI4.scala 171:24]
  assign io_out_arlock = 1'h0; // @[ToAXI4.scala 173:24]
  assign io_out_arcache = 4'h0; // @[ToAXI4.scala 174:24]
  assign io_out_arqos = 4'h0; // @[ToAXI4.scala 175:24]
  assign io_out_rready = io_in_resp_ready; // @[ToAXI4.scala 197:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  awAck = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wen = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      awAck <= 1'h0;
    end else if (wSend) begin
      awAck <= 1'h0;
    end else begin
      awAck <= _GEN_0;
    end
    if (reset) begin
      wAck <= 1'h0;
    end else if (wSend) begin
      wAck <= 1'h0;
    end else begin
      wAck <= _GEN_2;
    end
    if (_T_23) begin
      wen <= io_in_req_bits_cmd[0];
    end
  end
endmodule
module AXI4CLINT(
  input         clock,
  input         reset,
  output        io__in_awready,
  input         io__in_awvalid,
  input  [31:0] io__in_awaddr,
  output        io__in_wready,
  input         io__in_wvalid,
  input  [63:0] io__in_wdata,
  input  [7:0]  io__in_wstrb,
  input         io__in_bready,
  output        io__in_bvalid,
  output        io__in_arready,
  input         io__in_arvalid,
  input  [31:0] io__in_araddr,
  input         io__in_rready,
  output        io__in_rvalid,
  output [63:0] io__in_rdata,
  output        io__extra_mtip,
  output        io__extra_msip,
  output        io_extra_mtip,
  output        io_extra_msip
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [63:0] _RAND_5;
  reg [63:0] _RAND_6;
  reg [63:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
`endif // RANDOMIZE_REG_INIT
  wire [7:0] _T_9 = io__in_wstrb[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_11 = io__in_wstrb[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_13 = io__in_wstrb[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_15 = io__in_wstrb[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_17 = io__in_wstrb[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_19 = io__in_wstrb[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_21 = io__in_wstrb[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_23 = io__in_wstrb[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] fullMask = {_T_23,_T_21,_T_19,_T_17,_T_15,_T_13,_T_11,_T_9}; // @[Cat.scala 29:58]
  wire  _T_30 = io__in_arready & io__in_arvalid; // @[Decoupled.scala 40:37]
  wire  _T_31 = io__in_rready & io__in_rvalid; // @[Decoupled.scala 40:37]
  reg  r_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_31 ? 1'h0 : r_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_1 = _T_30 | _GEN_0; // @[StopWatch.scala 27:20]
  wire  _T_33 = ~r_busy; // @[AXI4Slave.scala 71:32]
  reg  ren; // @[AXI4Slave.scala 73:17]
  wire  _T_42 = _T_30 | r_busy; // @[AXI4Slave.scala 74:52]
  wire  _T_43 = ren & _T_42; // @[AXI4Slave.scala 74:35]
  reg  _T_45; // @[StopWatch.scala 24:20]
  wire  _GEN_2 = _T_31 ? 1'h0 : _T_45; // @[StopWatch.scala 26:19]
  wire  _GEN_3 = _T_43 | _GEN_2; // @[StopWatch.scala 27:20]
  wire  _T_46 = io__in_awready & io__in_awvalid; // @[Decoupled.scala 40:37]
  wire  _T_47 = io__in_bready & io__in_bvalid; // @[Decoupled.scala 40:37]
  reg  w_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_4 = _T_47 ? 1'h0 : w_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_5 = _T_46 | _GEN_4; // @[StopWatch.scala 27:20]
  wire  _T_50 = io__in_wready & io__in_wvalid; // @[Decoupled.scala 40:37]
  reg  _T_53; // @[StopWatch.scala 24:20]
  wire  _GEN_6 = _T_47 ? 1'h0 : _T_53; // @[StopWatch.scala 26:19]
  wire  _GEN_7 = _T_50 | _GEN_6; // @[StopWatch.scala 27:20]
  reg [63:0] mtime; // @[AXI4CLINT.scala 32:22]
  reg [63:0] mtimecmp; // @[AXI4CLINT.scala 33:25]
  reg [63:0] msip; // @[AXI4CLINT.scala 34:21]
  reg [15:0] freq; // @[AXI4CLINT.scala 37:21]
  reg [15:0] inc; // @[AXI4CLINT.scala 38:20]
  reg [15:0] cnt; // @[AXI4CLINT.scala 40:20]
  wire [15:0] nextCnt = cnt + 16'h1; // @[AXI4CLINT.scala 41:21]
  wire  _T_55 = nextCnt < freq; // @[AXI4CLINT.scala 42:22]
  wire  tick = nextCnt == freq; // @[AXI4CLINT.scala 43:23]
  wire [63:0] _GEN_14 = {{48'd0}, inc}; // @[AXI4CLINT.scala 44:32]
  wire [63:0] _T_58 = mtime + _GEN_14; // @[AXI4CLINT.scala 44:32]
  wire  _T_93 = 16'h0 == io__in_araddr[15:0]; // @[LookupTree.scala 24:34]
  wire  _T_94 = 16'h8000 == io__in_araddr[15:0]; // @[LookupTree.scala 24:34]
  wire  _T_95 = 16'hbff8 == io__in_araddr[15:0]; // @[LookupTree.scala 24:34]
  wire  _T_96 = 16'h8008 == io__in_araddr[15:0]; // @[LookupTree.scala 24:34]
  wire  _T_97 = 16'h4000 == io__in_araddr[15:0]; // @[LookupTree.scala 24:34]
  wire [63:0] _T_98 = _T_93 ? msip : 64'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_99 = _T_94 ? freq : 16'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_100 = _T_95 ? mtime : 64'h0; // @[Mux.scala 27:72]
  wire [15:0] _T_101 = _T_96 ? inc : 16'h0; // @[Mux.scala 27:72]
  wire [63:0] _T_102 = _T_97 ? mtimecmp : 64'h0; // @[Mux.scala 27:72]
  wire [63:0] _GEN_15 = {{48'd0}, _T_99}; // @[Mux.scala 27:72]
  wire [63:0] _T_103 = _T_98 | _GEN_15; // @[Mux.scala 27:72]
  wire [63:0] _T_104 = _T_103 | _T_100; // @[Mux.scala 27:72]
  wire [63:0] _GEN_16 = {{48'd0}, _T_101}; // @[Mux.scala 27:72]
  wire [63:0] _T_105 = _T_104 | _GEN_16; // @[Mux.scala 27:72]
  wire  _T_108 = io__in_awaddr[15:0] == 16'h0; // @[RegMap.scala 32:41]
  wire  _T_109 = _T_50 & _T_108; // @[RegMap.scala 32:32]
  wire [63:0] _T_110 = io__in_wdata & fullMask; // @[BitUtils.scala 32:13]
  wire [63:0] _T_111 = ~fullMask; // @[BitUtils.scala 32:38]
  wire [63:0] _T_112 = msip & _T_111; // @[BitUtils.scala 32:36]
  wire [63:0] _T_113 = _T_110 | _T_112; // @[BitUtils.scala 32:25]
  wire  _T_114 = io__in_awaddr[15:0] == 16'h8000; // @[RegMap.scala 32:41]
  wire  _T_115 = _T_50 & _T_114; // @[RegMap.scala 32:32]
  wire [63:0] _GEN_17 = {{48'd0}, freq}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_118 = _GEN_17 & _T_111; // @[BitUtils.scala 32:36]
  wire [63:0] _T_119 = _T_110 | _T_118; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_10 = _T_115 ? _T_119 : {{48'd0}, freq}; // @[RegMap.scala 32:48]
  wire  _T_120 = io__in_awaddr[15:0] == 16'hbff8; // @[RegMap.scala 32:41]
  wire  _T_121 = _T_50 & _T_120; // @[RegMap.scala 32:32]
  wire [63:0] _T_124 = mtime & _T_111; // @[BitUtils.scala 32:36]
  wire [63:0] _T_125 = _T_110 | _T_124; // @[BitUtils.scala 32:25]
  wire  _T_126 = io__in_awaddr[15:0] == 16'h8008; // @[RegMap.scala 32:41]
  wire  _T_127 = _T_50 & _T_126; // @[RegMap.scala 32:32]
  wire [63:0] _T_130 = _GEN_14 & _T_111; // @[BitUtils.scala 32:36]
  wire [63:0] _T_131 = _T_110 | _T_130; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_12 = _T_127 ? _T_131 : {{48'd0}, inc}; // @[RegMap.scala 32:48]
  wire  _T_132 = io__in_awaddr[15:0] == 16'h4000; // @[RegMap.scala 32:41]
  wire  _T_133 = _T_50 & _T_132; // @[RegMap.scala 32:32]
  wire [63:0] _T_136 = mtimecmp & _T_111; // @[BitUtils.scala 32:36]
  wire [63:0] _T_137 = _T_110 | _T_136; // @[BitUtils.scala 32:25]
  reg  _T_139; // @[AXI4CLINT.scala 64:31]
  reg  _T_141; // @[AXI4CLINT.scala 65:31]
  assign io__in_awready = ~w_busy; // @[AXI4Slave.scala 94:15]
  assign io__in_wready = io__in_awvalid | w_busy; // @[AXI4Slave.scala 95:15]
  assign io__in_bvalid = _T_53; // @[AXI4Slave.scala 97:14]
  assign io__in_arready = io__in_rready | _T_33; // @[AXI4Slave.scala 71:15]
  assign io__in_rvalid = _T_45; // @[AXI4Slave.scala 74:14]
  assign io__in_rdata = _T_105 | _T_102; // @[RegMap.scala 30:11]
  assign io__extra_mtip = _T_139; // @[AXI4CLINT.scala 64:21]
  assign io__extra_msip = _T_141; // @[AXI4CLINT.scala 65:21]
  assign io_extra_mtip = io__extra_mtip;
  assign io_extra_msip = io__extra_msip;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _T_45 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_53 = _RAND_4[0:0];
  _RAND_5 = {2{`RANDOM}};
  mtime = _RAND_5[63:0];
  _RAND_6 = {2{`RANDOM}};
  mtimecmp = _RAND_6[63:0];
  _RAND_7 = {2{`RANDOM}};
  msip = _RAND_7[63:0];
  _RAND_8 = {1{`RANDOM}};
  freq = _RAND_8[15:0];
  _RAND_9 = {1{`RANDOM}};
  inc = _RAND_9[15:0];
  _RAND_10 = {1{`RANDOM}};
  cnt = _RAND_10[15:0];
  _RAND_11 = {1{`RANDOM}};
  _T_139 = _RAND_11[0:0];
  _RAND_12 = {1{`RANDOM}};
  _T_141 = _RAND_12[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      r_busy <= 1'h0;
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin
      ren <= 1'h0;
    end else begin
      ren <= _T_30;
    end
    if (reset) begin
      _T_45 <= 1'h0;
    end else begin
      _T_45 <= _GEN_3;
    end
    if (reset) begin
      w_busy <= 1'h0;
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin
      _T_53 <= 1'h0;
    end else begin
      _T_53 <= _GEN_7;
    end
    if (reset) begin
      mtime <= 64'h0;
    end else if (_T_121) begin
      mtime <= _T_125;
    end else if (tick) begin
      mtime <= _T_58;
    end
    if (reset) begin
      mtimecmp <= 64'h0;
    end else if (_T_133) begin
      mtimecmp <= _T_137;
    end
    if (reset) begin
      msip <= 64'h0;
    end else if (_T_109) begin
      msip <= _T_113;
    end
    if (reset) begin
      freq <= 16'h28;
    end else begin
      freq <= _GEN_10[15:0];
    end
    if (reset) begin
      inc <= 16'h1;
    end else begin
      inc <= _GEN_12[15:0];
    end
    if (reset) begin
      cnt <= 16'h0;
    end else if (_T_55) begin
      cnt <= nextCnt;
    end else begin
      cnt <= 16'h0;
    end
    _T_139 <= mtime >= mtimecmp;
    _T_141 <= msip != 64'h0;
  end
endmodule
module SimpleBus2AXI4Converter_2(
  input         clock,
  input         reset,
  output        io_in_req_ready,
  input         io_in_req_valid,
  input  [31:0] io_in_req_bits_addr,
  input  [3:0]  io_in_req_bits_cmd,
  input  [7:0]  io_in_req_bits_wmask,
  input  [63:0] io_in_req_bits_wdata,
  input         io_in_resp_ready,
  output        io_in_resp_valid,
  output [63:0] io_in_resp_bits_rdata,
  input         io_out_awready,
  output        io_out_awvalid,
  output [31:0] io_out_awaddr,
  input         io_out_wready,
  output        io_out_wvalid,
  output [63:0] io_out_wdata,
  output [7:0]  io_out_wstrb,
  output        io_out_bready,
  input         io_out_bvalid,
  input         io_out_arready,
  output        io_out_arvalid,
  output [31:0] io_out_araddr,
  output        io_out_rready,
  input         io_out_rvalid,
  input  [63:0] io_out_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
`endif // RANDOMIZE_REG_INIT
  wire  _T_1 = io_in_req_valid & io_in_req_bits_cmd[1]; // @[ToAXI4.scala 151:38]
  wire  toAXI4Lite = ~_T_1; // @[ToAXI4.scala 151:20]
  wire  _T_5 = toAXI4Lite | reset; // @[ToAXI4.scala 153:9]
  wire  _T_6 = ~_T_5; // @[ToAXI4.scala 153:9]
  wire  _T_8 = io_out_awready & io_out_awvalid; // @[Decoupled.scala 40:37]
  reg  awAck; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_8 | awAck; // @[StopWatch.scala 30:20]
  wire  _T_12 = io_out_wready & io_out_wvalid; // @[Decoupled.scala 40:37]
  wire  _T_13 = _T_8 & _T_12; // @[ToAXI4.scala 189:27]
  reg  wAck; // @[StopWatch.scala 24:20]
  wire  _T_15 = awAck & wAck; // @[ToAXI4.scala 189:63]
  wire  wSend = _T_13 | _T_15; // @[ToAXI4.scala 189:53]
  wire  _GEN_2 = _T_12 | wAck; // @[StopWatch.scala 30:20]
  wire  _T_18 = io_in_req_ready & io_in_req_valid; // @[Decoupled.scala 40:37]
  reg  wen; // @[Reg.scala 15:16]
  wire  _T_20 = ~io_in_req_bits_cmd[0]; // @[SimpleBus.scala 73:18]
  wire  _T_22 = ~io_in_req_bits_cmd[3]; // @[SimpleBus.scala 73:29]
  wire  _T_23 = _T_20 & _T_22; // @[SimpleBus.scala 73:26]
  wire  _T_26 = io_in_req_valid & io_in_req_bits_cmd[0]; // @[SimpleBus.scala 103:29]
  wire  _T_27 = ~awAck; // @[ToAXI4.scala 193:36]
  wire  _T_31 = ~wAck; // @[ToAXI4.scala 194:36]
  wire  _T_35 = _T_31 & io_out_wready; // @[ToAXI4.scala 195:55]
  assign io_in_req_ready = io_in_req_bits_cmd[0] ? _T_35 : io_out_arready; // @[ToAXI4.scala 195:18]
  assign io_in_resp_valid = wen ? io_out_bvalid : io_out_rvalid; // @[ToAXI4.scala 199:19]
  assign io_in_resp_bits_rdata = io_out_rdata; // @[ToAXI4.scala 183:23]
  assign io_out_awvalid = _T_26 & _T_27; // @[ToAXI4.scala 193:16]
  assign io_out_awaddr = io_out_araddr; // @[ToAXI4.scala 182:6]
  assign io_out_wvalid = _T_26 & _T_31; // @[ToAXI4.scala 194:16]
  assign io_out_wdata = io_in_req_bits_wdata; // @[ToAXI4.scala 160:10]
  assign io_out_wstrb = io_in_req_bits_wmask; // @[ToAXI4.scala 161:10]
  assign io_out_bready = io_in_resp_ready; // @[ToAXI4.scala 198:16]
  assign io_out_arvalid = io_in_req_valid & _T_23; // @[ToAXI4.scala 192:16]
  assign io_out_araddr = io_in_req_bits_addr; // @[ToAXI4.scala 158:12]
  assign io_out_rready = io_in_resp_ready; // @[ToAXI4.scala 197:16]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  awAck = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  wAck = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  wen = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      awAck <= 1'h0;
    end else if (wSend) begin
      awAck <= 1'h0;
    end else begin
      awAck <= _GEN_0;
    end
    if (reset) begin
      wAck <= 1'h0;
    end else if (wSend) begin
      wAck <= 1'h0;
    end else begin
      wAck <= _GEN_2;
    end
    if (_T_18) begin
      wen <= io_in_req_bits_cmd[0];
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_6) begin
          $fwrite(32'h80000002,"Assertion failed\n    at ToAXI4.scala:153 assert(toAXI4Lite || toAXI4)\n"); // @[ToAXI4.scala 153:9]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_6) begin
          $fatal; // @[ToAXI4.scala 153:9]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module AXI4PLIC(
  input         clock,
  input         reset,
  output        io__in_awready,
  input         io__in_awvalid,
  input  [31:0] io__in_awaddr,
  output        io__in_wready,
  input         io__in_wvalid,
  input  [63:0] io__in_wdata,
  input  [7:0]  io__in_wstrb,
  input         io__in_bready,
  output        io__in_bvalid,
  output        io__in_arready,
  input         io__in_arvalid,
  input  [31:0] io__in_araddr,
  input         io__in_rready,
  output        io__in_rvalid,
  output [63:0] io__in_rdata,
  input  [2:0]  io__extra_intrVec,
  output        io__extra_meip_0,
  output        io_extra_meip_0
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_14;
  reg [31:0] _RAND_15;
  reg [31:0] _RAND_16;
`endif // RANDOMIZE_REG_INIT
  wire  _T_30 = io__in_arready & io__in_arvalid; // @[Decoupled.scala 40:37]
  wire  _T_31 = io__in_rready & io__in_rvalid; // @[Decoupled.scala 40:37]
  reg  r_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_31 ? 1'h0 : r_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_1 = _T_30 | _GEN_0; // @[StopWatch.scala 27:20]
  wire  _T_33 = ~r_busy; // @[AXI4Slave.scala 71:32]
  reg  ren; // @[AXI4Slave.scala 73:17]
  wire  _T_42 = _T_30 | r_busy; // @[AXI4Slave.scala 74:52]
  wire  _T_43 = ren & _T_42; // @[AXI4Slave.scala 74:35]
  reg  _T_45; // @[StopWatch.scala 24:20]
  wire  _GEN_2 = _T_31 ? 1'h0 : _T_45; // @[StopWatch.scala 26:19]
  wire  _GEN_3 = _T_43 | _GEN_2; // @[StopWatch.scala 27:20]
  wire  _T_46 = io__in_awready & io__in_awvalid; // @[Decoupled.scala 40:37]
  wire  _T_47 = io__in_bready & io__in_bvalid; // @[Decoupled.scala 40:37]
  reg  w_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_4 = _T_47 ? 1'h0 : w_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_5 = _T_46 | _GEN_4; // @[StopWatch.scala 27:20]
  wire  _T_50 = io__in_wready & io__in_wvalid; // @[Decoupled.scala 40:37]
  reg  _T_53; // @[StopWatch.scala 24:20]
  wire  _GEN_6 = _T_47 ? 1'h0 : _T_53; // @[StopWatch.scala 26:19]
  wire  _GEN_7 = _T_50 | _GEN_6; // @[StopWatch.scala 27:20]
  reg [31:0] priority_0; // @[AXI4PLIC.scala 37:39]
  reg [31:0] priority_1; // @[AXI4PLIC.scala 37:39]
  reg [31:0] priority_2; // @[AXI4PLIC.scala 37:39]
  reg  pending_0_1; // @[AXI4PLIC.scala 43:46]
  reg  pending_0_2; // @[AXI4PLIC.scala 43:46]
  reg  pending_0_3; // @[AXI4PLIC.scala 43:46]
  wire [31:0] _T_85 = {16'h0,8'h0,4'h0,pending_0_3,pending_0_2,pending_0_1,1'h0}; // @[Cat.scala 29:58]
  reg [31:0] enable_0_0; // @[AXI4PLIC.scala 48:64]
  reg [31:0] threshold_0; // @[AXI4PLIC.scala 53:40]
  reg  inHandle_1; // @[AXI4PLIC.scala 58:25]
  reg  inHandle_2; // @[AXI4PLIC.scala 58:25]
  reg  inHandle_3; // @[AXI4PLIC.scala 58:25]
  reg [31:0] claimCompletion_0; // @[AXI4PLIC.scala 64:46]
  wire  _T_89 = io__in_araddr[25:0] == 26'h200004; // @[AXI4PLIC.scala 68:46]
  wire  _T_90 = _T_31 & _T_89; // @[AXI4PLIC.scala 68:25]
  wire  _GEN_37 = 2'h1 == claimCompletion_0[1:0]; // @[AXI4PLIC.scala 68:73]
  wire  _GEN_9 = _GEN_37 | inHandle_1; // @[AXI4PLIC.scala 68:73]
  wire  _GEN_38 = 2'h2 == claimCompletion_0[1:0]; // @[AXI4PLIC.scala 68:73]
  wire  _GEN_10 = _GEN_38 | inHandle_2; // @[AXI4PLIC.scala 68:73]
  wire  _GEN_39 = 2'h3 == claimCompletion_0[1:0]; // @[AXI4PLIC.scala 68:73]
  wire  _GEN_11 = _GEN_39 | inHandle_3; // @[AXI4PLIC.scala 68:73]
  wire  _GEN_16 = io__extra_intrVec[0] | pending_0_1; // @[AXI4PLIC.scala 75:17]
  wire  _GEN_18 = io__extra_intrVec[1] | pending_0_2; // @[AXI4PLIC.scala 75:17]
  wire  _GEN_20 = io__extra_intrVec[2] | pending_0_3; // @[AXI4PLIC.scala 75:17]
  wire [31:0] _T_125 = _T_85 & enable_0_0; // @[AXI4PLIC.scala 81:31]
  wire  _T_126 = _T_125 == 32'h0; // @[AXI4PLIC.scala 82:23]
  wire [4:0] _T_159 = _T_125[30] ? 5'h1e : 5'h1f; // @[Mux.scala 47:69]
  wire [4:0] _T_160 = _T_125[29] ? 5'h1d : _T_159; // @[Mux.scala 47:69]
  wire [4:0] _T_161 = _T_125[28] ? 5'h1c : _T_160; // @[Mux.scala 47:69]
  wire [4:0] _T_162 = _T_125[27] ? 5'h1b : _T_161; // @[Mux.scala 47:69]
  wire [4:0] _T_163 = _T_125[26] ? 5'h1a : _T_162; // @[Mux.scala 47:69]
  wire [4:0] _T_164 = _T_125[25] ? 5'h19 : _T_163; // @[Mux.scala 47:69]
  wire [4:0] _T_165 = _T_125[24] ? 5'h18 : _T_164; // @[Mux.scala 47:69]
  wire [4:0] _T_166 = _T_125[23] ? 5'h17 : _T_165; // @[Mux.scala 47:69]
  wire [4:0] _T_167 = _T_125[22] ? 5'h16 : _T_166; // @[Mux.scala 47:69]
  wire [4:0] _T_168 = _T_125[21] ? 5'h15 : _T_167; // @[Mux.scala 47:69]
  wire [4:0] _T_169 = _T_125[20] ? 5'h14 : _T_168; // @[Mux.scala 47:69]
  wire [4:0] _T_170 = _T_125[19] ? 5'h13 : _T_169; // @[Mux.scala 47:69]
  wire [4:0] _T_171 = _T_125[18] ? 5'h12 : _T_170; // @[Mux.scala 47:69]
  wire [4:0] _T_172 = _T_125[17] ? 5'h11 : _T_171; // @[Mux.scala 47:69]
  wire [4:0] _T_173 = _T_125[16] ? 5'h10 : _T_172; // @[Mux.scala 47:69]
  wire [4:0] _T_174 = _T_125[15] ? 5'hf : _T_173; // @[Mux.scala 47:69]
  wire [4:0] _T_175 = _T_125[14] ? 5'he : _T_174; // @[Mux.scala 47:69]
  wire [4:0] _T_176 = _T_125[13] ? 5'hd : _T_175; // @[Mux.scala 47:69]
  wire [4:0] _T_177 = _T_125[12] ? 5'hc : _T_176; // @[Mux.scala 47:69]
  wire [4:0] _T_178 = _T_125[11] ? 5'hb : _T_177; // @[Mux.scala 47:69]
  wire [4:0] _T_179 = _T_125[10] ? 5'ha : _T_178; // @[Mux.scala 47:69]
  wire [4:0] _T_180 = _T_125[9] ? 5'h9 : _T_179; // @[Mux.scala 47:69]
  wire [4:0] _T_181 = _T_125[8] ? 5'h8 : _T_180; // @[Mux.scala 47:69]
  wire [4:0] _T_182 = _T_125[7] ? 5'h7 : _T_181; // @[Mux.scala 47:69]
  wire [4:0] _T_183 = _T_125[6] ? 5'h6 : _T_182; // @[Mux.scala 47:69]
  wire [4:0] _T_184 = _T_125[5] ? 5'h5 : _T_183; // @[Mux.scala 47:69]
  wire [4:0] _T_185 = _T_125[4] ? 5'h4 : _T_184; // @[Mux.scala 47:69]
  wire [4:0] _T_186 = _T_125[3] ? 5'h3 : _T_185; // @[Mux.scala 47:69]
  wire [4:0] _T_187 = _T_125[2] ? 5'h2 : _T_186; // @[Mux.scala 47:69]
  wire [4:0] _T_188 = _T_125[1] ? 5'h1 : _T_187; // @[Mux.scala 47:69]
  wire [4:0] _T_189 = _T_125[0] ? 5'h0 : _T_188; // @[Mux.scala 47:69]
  wire [4:0] _T_190 = _T_126 ? 5'h0 : _T_189; // @[AXI4PLIC.scala 82:13]
  wire [7:0] _T_195 = io__in_wstrb >> io__in_awaddr[2:0]; // @[AXI4PLIC.scala 89:78]
  wire [7:0] _T_205 = _T_195[0] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_207 = _T_195[1] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_209 = _T_195[2] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_211 = _T_195[3] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_213 = _T_195[4] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_215 = _T_195[5] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_217 = _T_195[6] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [7:0] _T_219 = _T_195[7] ? 8'hff : 8'h0; // @[Bitwise.scala 72:12]
  wire [63:0] _T_226 = {_T_219,_T_217,_T_215,_T_213,_T_211,_T_209,_T_207,_T_205}; // @[Cat.scala 29:58]
  wire  _T_227 = 26'hc == io__in_araddr[25:0]; // @[LookupTree.scala 24:34]
  wire  _T_228 = 26'h1000 == io__in_araddr[25:0]; // @[LookupTree.scala 24:34]
  wire  _T_229 = 26'h2000 == io__in_araddr[25:0]; // @[LookupTree.scala 24:34]
  wire  _T_230 = 26'h8 == io__in_araddr[25:0]; // @[LookupTree.scala 24:34]
  wire  _T_231 = 26'h200004 == io__in_araddr[25:0]; // @[LookupTree.scala 24:34]
  wire  _T_232 = 26'h4 == io__in_araddr[25:0]; // @[LookupTree.scala 24:34]
  wire  _T_233 = 26'h200000 == io__in_araddr[25:0]; // @[LookupTree.scala 24:34]
  wire [31:0] _T_234 = _T_227 ? priority_2 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_235 = _T_228 ? _T_85 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_236 = _T_229 ? enable_0_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_237 = _T_230 ? priority_1 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_238 = _T_231 ? claimCompletion_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_239 = _T_232 ? priority_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_240 = _T_233 ? threshold_0 : 32'h0; // @[Mux.scala 27:72]
  wire [31:0] _T_241 = _T_234 | _T_235; // @[Mux.scala 27:72]
  wire [31:0] _T_242 = _T_241 | _T_236; // @[Mux.scala 27:72]
  wire [31:0] _T_243 = _T_242 | _T_237; // @[Mux.scala 27:72]
  wire [31:0] _T_244 = _T_243 | _T_238; // @[Mux.scala 27:72]
  wire [31:0] _T_245 = _T_244 | _T_239; // @[Mux.scala 27:72]
  wire [31:0] rdata = _T_245 | _T_240; // @[Mux.scala 27:72]
  wire  _T_248 = io__in_awaddr[25:0] == 26'hc; // @[RegMap.scala 32:41]
  wire  _T_249 = _T_50 & _T_248; // @[RegMap.scala 32:32]
  wire [63:0] _T_250 = io__in_wdata & _T_226; // @[BitUtils.scala 32:13]
  wire [63:0] _T_251 = ~_T_226; // @[BitUtils.scala 32:38]
  wire [63:0] _GEN_40 = {{32'd0}, priority_2}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_252 = _GEN_40 & _T_251; // @[BitUtils.scala 32:36]
  wire [63:0] _T_253 = _T_250 | _T_252; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_22 = _T_249 ? _T_253 : {{32'd0}, priority_2}; // @[RegMap.scala 32:48]
  wire  _T_254 = io__in_awaddr[25:0] == 26'h2000; // @[RegMap.scala 32:41]
  wire  _T_255 = _T_50 & _T_254; // @[RegMap.scala 32:32]
  wire [63:0] _GEN_41 = {{32'd0}, enable_0_0}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_258 = _GEN_41 & _T_251; // @[BitUtils.scala 32:36]
  wire [63:0] _T_259 = _T_250 | _T_258; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_23 = _T_255 ? _T_259 : {{32'd0}, enable_0_0}; // @[RegMap.scala 32:48]
  wire  _T_260 = io__in_awaddr[25:0] == 26'h8; // @[RegMap.scala 32:41]
  wire  _T_261 = _T_50 & _T_260; // @[RegMap.scala 32:32]
  wire [63:0] _GEN_42 = {{32'd0}, priority_1}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_264 = _GEN_42 & _T_251; // @[BitUtils.scala 32:36]
  wire [63:0] _T_265 = _T_250 | _T_264; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_24 = _T_261 ? _T_265 : {{32'd0}, priority_1}; // @[RegMap.scala 32:48]
  wire  _T_266 = io__in_awaddr[25:0] == 26'h200004; // @[RegMap.scala 32:41]
  wire  _T_267 = _T_50 & _T_266; // @[RegMap.scala 32:32]
  wire [63:0] _GEN_43 = {{32'd0}, claimCompletion_0}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_270 = _GEN_43 & _T_251; // @[BitUtils.scala 32:36]
  wire [63:0] _T_271 = _T_250 | _T_270; // @[BitUtils.scala 32:25]
  wire [4:0] _GEN_33 = _T_267 ? 5'h0 : _T_190; // @[RegMap.scala 32:48]
  wire  _T_274 = io__in_awaddr[25:0] == 26'h4; // @[RegMap.scala 32:41]
  wire  _T_275 = _T_50 & _T_274; // @[RegMap.scala 32:32]
  wire [63:0] _GEN_44 = {{32'd0}, priority_0}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_278 = _GEN_44 & _T_251; // @[BitUtils.scala 32:36]
  wire [63:0] _T_279 = _T_250 | _T_278; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_34 = _T_275 ? _T_279 : {{32'd0}, priority_0}; // @[RegMap.scala 32:48]
  wire  _T_280 = io__in_awaddr[25:0] == 26'h200000; // @[RegMap.scala 32:41]
  wire  _T_281 = _T_50 & _T_280; // @[RegMap.scala 32:32]
  wire [63:0] _GEN_45 = {{32'd0}, threshold_0}; // @[BitUtils.scala 32:36]
  wire [63:0] _T_284 = _GEN_45 & _T_251; // @[BitUtils.scala 32:36]
  wire [63:0] _T_285 = _T_250 | _T_284; // @[BitUtils.scala 32:25]
  wire [63:0] _GEN_35 = _T_281 ? _T_285 : {{32'd0}, threshold_0}; // @[RegMap.scala 32:48]
  assign io__in_awready = ~w_busy; // @[AXI4Slave.scala 94:15]
  assign io__in_wready = io__in_awvalid | w_busy; // @[AXI4Slave.scala 95:15]
  assign io__in_bvalid = _T_53; // @[AXI4Slave.scala 97:14]
  assign io__in_arready = io__in_rready | _T_33; // @[AXI4Slave.scala 71:15]
  assign io__in_rvalid = _T_45; // @[AXI4Slave.scala 74:14]
  assign io__in_rdata = {rdata,rdata}; // @[AXI4PLIC.scala 91:18]
  assign io__extra_meip_0 = claimCompletion_0 != 32'h0; // @[AXI4PLIC.scala 93:62]
  assign io_extra_meip_0 = io__extra_meip_0;
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _T_45 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_53 = _RAND_4[0:0];
  _RAND_5 = {1{`RANDOM}};
  priority_0 = _RAND_5[31:0];
  _RAND_6 = {1{`RANDOM}};
  priority_1 = _RAND_6[31:0];
  _RAND_7 = {1{`RANDOM}};
  priority_2 = _RAND_7[31:0];
  _RAND_8 = {1{`RANDOM}};
  pending_0_1 = _RAND_8[0:0];
  _RAND_9 = {1{`RANDOM}};
  pending_0_2 = _RAND_9[0:0];
  _RAND_10 = {1{`RANDOM}};
  pending_0_3 = _RAND_10[0:0];
  _RAND_11 = {1{`RANDOM}};
  enable_0_0 = _RAND_11[31:0];
  _RAND_12 = {1{`RANDOM}};
  threshold_0 = _RAND_12[31:0];
  _RAND_13 = {1{`RANDOM}};
  inHandle_1 = _RAND_13[0:0];
  _RAND_14 = {1{`RANDOM}};
  inHandle_2 = _RAND_14[0:0];
  _RAND_15 = {1{`RANDOM}};
  inHandle_3 = _RAND_15[0:0];
  _RAND_16 = {1{`RANDOM}};
  claimCompletion_0 = _RAND_16[31:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      r_busy <= 1'h0;
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin
      ren <= 1'h0;
    end else begin
      ren <= _T_30;
    end
    if (reset) begin
      _T_45 <= 1'h0;
    end else begin
      _T_45 <= _GEN_3;
    end
    if (reset) begin
      w_busy <= 1'h0;
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin
      _T_53 <= 1'h0;
    end else begin
      _T_53 <= _GEN_7;
    end
    priority_0 <= _GEN_34[31:0];
    priority_1 <= _GEN_24[31:0];
    priority_2 <= _GEN_22[31:0];
    if (reset) begin
      pending_0_1 <= 1'h0;
    end else if (inHandle_1) begin
      pending_0_1 <= 1'h0;
    end else begin
      pending_0_1 <= _GEN_16;
    end
    if (reset) begin
      pending_0_2 <= 1'h0;
    end else if (inHandle_2) begin
      pending_0_2 <= 1'h0;
    end else begin
      pending_0_2 <= _GEN_18;
    end
    if (reset) begin
      pending_0_3 <= 1'h0;
    end else if (inHandle_3) begin
      pending_0_3 <= 1'h0;
    end else begin
      pending_0_3 <= _GEN_20;
    end
    if (reset) begin
      enable_0_0 <= 32'h0;
    end else begin
      enable_0_0 <= _GEN_23[31:0];
    end
    threshold_0 <= _GEN_35[31:0];
    if (reset) begin
      inHandle_1 <= 1'h0;
    end else if (_T_267) begin
      if (2'h1 == _T_271[1:0]) begin
        inHandle_1 <= 1'h0;
      end else if (_T_90) begin
        inHandle_1 <= _GEN_9;
      end
    end else if (_T_90) begin
      inHandle_1 <= _GEN_9;
    end
    if (reset) begin
      inHandle_2 <= 1'h0;
    end else if (_T_267) begin
      if (2'h2 == _T_271[1:0]) begin
        inHandle_2 <= 1'h0;
      end else if (_T_90) begin
        inHandle_2 <= _GEN_10;
      end
    end else if (_T_90) begin
      inHandle_2 <= _GEN_10;
    end
    if (reset) begin
      inHandle_3 <= 1'h0;
    end else if (_T_267) begin
      if (2'h3 == _T_271[1:0]) begin
        inHandle_3 <= 1'h0;
      end else if (_T_90) begin
        inHandle_3 <= _GEN_11;
      end
    end else if (_T_90) begin
      inHandle_3 <= _GEN_11;
    end
    claimCompletion_0 <= {{27'd0}, _GEN_33};
  end
endmodule
module NutShell(
  input         clock,
  input         reset,
  input         io_mem_awready,
  output        io_mem_awvalid,
  output [31:0] io_mem_awaddr,
  output [2:0]  io_mem_awprot,
  output        io_mem_awid,
  output        io_mem_awuser,
  output [7:0]  io_mem_awlen,
  output [2:0]  io_mem_awsize,
  output [1:0]  io_mem_awburst,
  output        io_mem_awlock,
  output [3:0]  io_mem_awcache,
  output [3:0]  io_mem_awqos,
  input         io_mem_wready,
  output        io_mem_wvalid,
  output [63:0] io_mem_wdata,
  output [7:0]  io_mem_wstrb,
  output        io_mem_wlast,
  output        io_mem_bready,
  input         io_mem_bvalid,
  input  [1:0]  io_mem_bresp,
  input         io_mem_bid,
  input         io_mem_buser,
  input         io_mem_arready,
  output        io_mem_arvalid,
  output [31:0] io_mem_araddr,
  output [2:0]  io_mem_arprot,
  output        io_mem_arid,
  output        io_mem_aruser,
  output [7:0]  io_mem_arlen,
  output [2:0]  io_mem_arsize,
  output [1:0]  io_mem_arburst,
  output        io_mem_arlock,
  output [3:0]  io_mem_arcache,
  output [3:0]  io_mem_arqos,
  output        io_mem_rready,
  input         io_mem_rvalid,
  input  [1:0]  io_mem_rresp,
  input  [63:0] io_mem_rdata,
  input         io_mem_rlast,
  input         io_mem_rid,
  input         io_mem_ruser,
  input         io_mmio_awready,
  output        io_mmio_awvalid,
  output [31:0] io_mmio_awaddr,
  output [2:0]  io_mmio_awprot,
  output        io_mmio_awid,
  output        io_mmio_awuser,
  output [7:0]  io_mmio_awlen,
  output [2:0]  io_mmio_awsize,
  output [1:0]  io_mmio_awburst,
  output        io_mmio_awlock,
  output [3:0]  io_mmio_awcache,
  output [3:0]  io_mmio_awqos,
  input         io_mmio_wready,
  output        io_mmio_wvalid,
  output [63:0] io_mmio_wdata,
  output [7:0]  io_mmio_wstrb,
  output        io_mmio_wlast,
  output        io_mmio_bready,
  input         io_mmio_bvalid,
  input  [1:0]  io_mmio_bresp,
  input         io_mmio_bid,
  input         io_mmio_buser,
  input         io_mmio_arready,
  output        io_mmio_arvalid,
  output [31:0] io_mmio_araddr,
  output [2:0]  io_mmio_arprot,
  output        io_mmio_arid,
  output        io_mmio_aruser,
  output [7:0]  io_mmio_arlen,
  output [2:0]  io_mmio_arsize,
  output [1:0]  io_mmio_arburst,
  output        io_mmio_arlock,
  output [3:0]  io_mmio_arcache,
  output [3:0]  io_mmio_arqos,
  output        io_mmio_rready,
  input         io_mmio_rvalid,
  input  [1:0]  io_mmio_rresp,
  input  [63:0] io_mmio_rdata,
  input         io_mmio_rlast,
  input         io_mmio_rid,
  input         io_mmio_ruser,
  output        io_frontend_awready,
  input         io_frontend_awvalid,
  input  [31:0] io_frontend_awaddr,
  input  [2:0]  io_frontend_awprot,
  input         io_frontend_awid,
  input         io_frontend_awuser,
  input  [7:0]  io_frontend_awlen,
  input  [2:0]  io_frontend_awsize,
  input  [1:0]  io_frontend_awburst,
  input         io_frontend_awlock,
  input  [3:0]  io_frontend_awcache,
  input  [3:0]  io_frontend_awqos,
  output        io_frontend_wready,
  input         io_frontend_wvalid,
  input  [63:0] io_frontend_wdata,
  input  [7:0]  io_frontend_wstrb,
  input         io_frontend_wlast,
  input         io_frontend_bready,
  output        io_frontend_bvalid,
  output [1:0]  io_frontend_bresp,
  output        io_frontend_bid,
  output        io_frontend_buser,
  output        io_frontend_arready,
  input         io_frontend_arvalid,
  input  [31:0] io_frontend_araddr,
  input  [2:0]  io_frontend_arprot,
  input         io_frontend_arid,
  input         io_frontend_aruser,
  input  [7:0]  io_frontend_arlen,
  input  [2:0]  io_frontend_arsize,
  input  [1:0]  io_frontend_arburst,
  input         io_frontend_arlock,
  input  [3:0]  io_frontend_arcache,
  input  [3:0]  io_frontend_arqos,
  input         io_frontend_rready,
  output        io_frontend_rvalid,
  output [1:0]  io_frontend_rresp,
  output [63:0] io_frontend_rdata,
  output        io_frontend_rlast,
  output        io_frontend_rid,
  output        io_frontend_ruser,
  input  [2:0]  io_meip,
  output [38:0] io_ila_WBUpc,
  output        io_ila_WBUvalid,
  output        io_ila_WBUrfWen,
  output [4:0]  io_ila_WBUrfDest,
  output [63:0] io_ila_WBUrfData,
  output [63:0] io_ila_InstrCnt
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
`endif // RANDOMIZE_REG_INIT
  wire  nutcore_clock; // @[NutShell.scala 53:23]
  wire  nutcore_reset; // @[NutShell.scala 53:23]
  wire  nutcore_io_imem_mem_req_ready; // @[NutShell.scala 53:23]
  wire  nutcore_io_imem_mem_req_valid; // @[NutShell.scala 53:23]
  wire [31:0] nutcore_io_imem_mem_req_bits_addr; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_imem_mem_req_bits_cmd; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_imem_mem_req_bits_wdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_imem_mem_resp_valid; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_imem_mem_resp_bits_cmd; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_imem_mem_resp_bits_rdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_dmem_mem_req_ready; // @[NutShell.scala 53:23]
  wire  nutcore_io_dmem_mem_req_valid; // @[NutShell.scala 53:23]
  wire [31:0] nutcore_io_dmem_mem_req_bits_addr; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_dmem_mem_req_bits_cmd; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_dmem_mem_req_bits_wdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_dmem_mem_resp_valid; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_dmem_mem_resp_bits_cmd; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_dmem_mem_resp_bits_rdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_dmem_coh_req_ready; // @[NutShell.scala 53:23]
  wire  nutcore_io_dmem_coh_req_valid; // @[NutShell.scala 53:23]
  wire [31:0] nutcore_io_dmem_coh_req_bits_addr; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_dmem_coh_req_bits_wdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_dmem_coh_resp_valid; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_dmem_coh_resp_bits_cmd; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_dmem_coh_resp_bits_rdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_mmio_req_ready; // @[NutShell.scala 53:23]
  wire  nutcore_io_mmio_req_valid; // @[NutShell.scala 53:23]
  wire [31:0] nutcore_io_mmio_req_bits_addr; // @[NutShell.scala 53:23]
  wire [2:0] nutcore_io_mmio_req_bits_size; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_mmio_req_bits_cmd; // @[NutShell.scala 53:23]
  wire [7:0] nutcore_io_mmio_req_bits_wmask; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_mmio_req_bits_wdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_mmio_resp_valid; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_mmio_resp_bits_cmd; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_mmio_resp_bits_rdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_frontend_req_ready; // @[NutShell.scala 53:23]
  wire  nutcore_io_frontend_req_valid; // @[NutShell.scala 53:23]
  wire [31:0] nutcore_io_frontend_req_bits_addr; // @[NutShell.scala 53:23]
  wire [2:0] nutcore_io_frontend_req_bits_size; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_frontend_req_bits_cmd; // @[NutShell.scala 53:23]
  wire [7:0] nutcore_io_frontend_req_bits_wmask; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_frontend_req_bits_wdata; // @[NutShell.scala 53:23]
  wire  nutcore_io_frontend_resp_ready; // @[NutShell.scala 53:23]
  wire  nutcore_io_frontend_resp_valid; // @[NutShell.scala 53:23]
  wire [3:0] nutcore_io_frontend_resp_bits_cmd; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_frontend_resp_bits_rdata; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_perfCnts_2; // @[NutShell.scala 53:23]
  wire [38:0] nutcore_io_in_bits_decode_cf_pc; // @[NutShell.scala 53:23]
  wire [4:0] nutcore_io_wb_rfDest; // @[NutShell.scala 53:23]
  wire  nutcore_io_extra_mtip; // @[NutShell.scala 53:23]
  wire  nutcore_io_extra_meip_0; // @[NutShell.scala 53:23]
  wire  nutcore_io_wb_rfWen; // @[NutShell.scala 53:23]
  wire [63:0] nutcore_io_wb_rfData; // @[NutShell.scala 53:23]
  wire  nutcore_io_extra_msip; // @[NutShell.scala 53:23]
  wire  nutcore_io_in_valid_0; // @[NutShell.scala 53:23]
  wire  cohMg_clock; // @[NutShell.scala 54:21]
  wire  cohMg_reset; // @[NutShell.scala 54:21]
  wire  cohMg_io_in_req_ready; // @[NutShell.scala 54:21]
  wire  cohMg_io_in_req_valid; // @[NutShell.scala 54:21]
  wire [31:0] cohMg_io_in_req_bits_addr; // @[NutShell.scala 54:21]
  wire [3:0] cohMg_io_in_req_bits_cmd; // @[NutShell.scala 54:21]
  wire [63:0] cohMg_io_in_req_bits_wdata; // @[NutShell.scala 54:21]
  wire  cohMg_io_in_resp_valid; // @[NutShell.scala 54:21]
  wire [3:0] cohMg_io_in_resp_bits_cmd; // @[NutShell.scala 54:21]
  wire [63:0] cohMg_io_in_resp_bits_rdata; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_mem_req_ready; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_mem_req_valid; // @[NutShell.scala 54:21]
  wire [31:0] cohMg_io_out_mem_req_bits_addr; // @[NutShell.scala 54:21]
  wire [3:0] cohMg_io_out_mem_req_bits_cmd; // @[NutShell.scala 54:21]
  wire [63:0] cohMg_io_out_mem_req_bits_wdata; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_mem_resp_ready; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_mem_resp_valid; // @[NutShell.scala 54:21]
  wire [3:0] cohMg_io_out_mem_resp_bits_cmd; // @[NutShell.scala 54:21]
  wire [63:0] cohMg_io_out_mem_resp_bits_rdata; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_coh_req_ready; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_coh_req_valid; // @[NutShell.scala 54:21]
  wire [31:0] cohMg_io_out_coh_req_bits_addr; // @[NutShell.scala 54:21]
  wire [63:0] cohMg_io_out_coh_req_bits_wdata; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_coh_resp_ready; // @[NutShell.scala 54:21]
  wire  cohMg_io_out_coh_resp_valid; // @[NutShell.scala 54:21]
  wire [3:0] cohMg_io_out_coh_resp_bits_cmd; // @[NutShell.scala 54:21]
  wire [63:0] cohMg_io_out_coh_resp_bits_rdata; // @[NutShell.scala 54:21]
  wire  xbar_clock; // @[NutShell.scala 55:20]
  wire  xbar_reset; // @[NutShell.scala 55:20]
  wire  xbar_io_in_0_req_ready; // @[NutShell.scala 55:20]
  wire  xbar_io_in_0_req_valid; // @[NutShell.scala 55:20]
  wire [31:0] xbar_io_in_0_req_bits_addr; // @[NutShell.scala 55:20]
  wire [3:0] xbar_io_in_0_req_bits_cmd; // @[NutShell.scala 55:20]
  wire [7:0] xbar_io_in_0_req_bits_wmask; // @[NutShell.scala 55:20]
  wire [63:0] xbar_io_in_0_req_bits_wdata; // @[NutShell.scala 55:20]
  wire  xbar_io_in_0_resp_valid; // @[NutShell.scala 55:20]
  wire [3:0] xbar_io_in_0_resp_bits_cmd; // @[NutShell.scala 55:20]
  wire [63:0] xbar_io_in_0_resp_bits_rdata; // @[NutShell.scala 55:20]
  wire  xbar_io_in_1_req_ready; // @[NutShell.scala 55:20]
  wire  xbar_io_in_1_req_valid; // @[NutShell.scala 55:20]
  wire [31:0] xbar_io_in_1_req_bits_addr; // @[NutShell.scala 55:20]
  wire [2:0] xbar_io_in_1_req_bits_size; // @[NutShell.scala 55:20]
  wire [3:0] xbar_io_in_1_req_bits_cmd; // @[NutShell.scala 55:20]
  wire [7:0] xbar_io_in_1_req_bits_wmask; // @[NutShell.scala 55:20]
  wire [63:0] xbar_io_in_1_req_bits_wdata; // @[NutShell.scala 55:20]
  wire  xbar_io_in_1_resp_valid; // @[NutShell.scala 55:20]
  wire [3:0] xbar_io_in_1_resp_bits_cmd; // @[NutShell.scala 55:20]
  wire [63:0] xbar_io_in_1_resp_bits_rdata; // @[NutShell.scala 55:20]
  wire  xbar_io_out_req_ready; // @[NutShell.scala 55:20]
  wire  xbar_io_out_req_valid; // @[NutShell.scala 55:20]
  wire [31:0] xbar_io_out_req_bits_addr; // @[NutShell.scala 55:20]
  wire [2:0] xbar_io_out_req_bits_size; // @[NutShell.scala 55:20]
  wire [3:0] xbar_io_out_req_bits_cmd; // @[NutShell.scala 55:20]
  wire [7:0] xbar_io_out_req_bits_wmask; // @[NutShell.scala 55:20]
  wire [63:0] xbar_io_out_req_bits_wdata; // @[NutShell.scala 55:20]
  wire  xbar_io_out_resp_ready; // @[NutShell.scala 55:20]
  wire  xbar_io_out_resp_valid; // @[NutShell.scala 55:20]
  wire [3:0] xbar_io_out_resp_bits_cmd; // @[NutShell.scala 55:20]
  wire [63:0] xbar_io_out_resp_bits_rdata; // @[NutShell.scala 55:20]
  wire  axi2sb_clock; // @[NutShell.scala 61:22]
  wire  axi2sb_reset; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_awready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_awvalid; // @[NutShell.scala 61:22]
  wire [31:0] axi2sb_io_in_awaddr; // @[NutShell.scala 61:22]
  wire [17:0] axi2sb_io_in_awid; // @[NutShell.scala 61:22]
  wire [7:0] axi2sb_io_in_awlen; // @[NutShell.scala 61:22]
  wire [2:0] axi2sb_io_in_awsize; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_wready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_wvalid; // @[NutShell.scala 61:22]
  wire [63:0] axi2sb_io_in_wdata; // @[NutShell.scala 61:22]
  wire [7:0] axi2sb_io_in_wstrb; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_wlast; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_bready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_bvalid; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_arready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_arvalid; // @[NutShell.scala 61:22]
  wire [31:0] axi2sb_io_in_araddr; // @[NutShell.scala 61:22]
  wire [17:0] axi2sb_io_in_arid; // @[NutShell.scala 61:22]
  wire [7:0] axi2sb_io_in_arlen; // @[NutShell.scala 61:22]
  wire [2:0] axi2sb_io_in_arsize; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_rready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_rvalid; // @[NutShell.scala 61:22]
  wire [63:0] axi2sb_io_in_rdata; // @[NutShell.scala 61:22]
  wire  axi2sb_io_in_rlast; // @[NutShell.scala 61:22]
  wire [17:0] axi2sb_io_in_rid; // @[NutShell.scala 61:22]
  wire  axi2sb_io_out_req_ready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_out_req_valid; // @[NutShell.scala 61:22]
  wire [31:0] axi2sb_io_out_req_bits_addr; // @[NutShell.scala 61:22]
  wire [2:0] axi2sb_io_out_req_bits_size; // @[NutShell.scala 61:22]
  wire [3:0] axi2sb_io_out_req_bits_cmd; // @[NutShell.scala 61:22]
  wire [7:0] axi2sb_io_out_req_bits_wmask; // @[NutShell.scala 61:22]
  wire [63:0] axi2sb_io_out_req_bits_wdata; // @[NutShell.scala 61:22]
  wire  axi2sb_io_out_resp_ready; // @[NutShell.scala 61:22]
  wire  axi2sb_io_out_resp_valid; // @[NutShell.scala 61:22]
  wire [3:0] axi2sb_io_out_resp_bits_cmd; // @[NutShell.scala 61:22]
  wire [63:0] axi2sb_io_out_resp_bits_rdata; // @[NutShell.scala 61:22]
  wire  Prefetcher_clock; // @[NutShell.scala 73:30]
  wire  Prefetcher_reset; // @[NutShell.scala 73:30]
  wire  Prefetcher_io_in_ready; // @[NutShell.scala 73:30]
  wire  Prefetcher_io_in_valid; // @[NutShell.scala 73:30]
  wire [31:0] Prefetcher_io_in_bits_addr; // @[NutShell.scala 73:30]
  wire [2:0] Prefetcher_io_in_bits_size; // @[NutShell.scala 73:30]
  wire [3:0] Prefetcher_io_in_bits_cmd; // @[NutShell.scala 73:30]
  wire [7:0] Prefetcher_io_in_bits_wmask; // @[NutShell.scala 73:30]
  wire [63:0] Prefetcher_io_in_bits_wdata; // @[NutShell.scala 73:30]
  wire  Prefetcher_io_out_ready; // @[NutShell.scala 73:30]
  wire  Prefetcher_io_out_valid; // @[NutShell.scala 73:30]
  wire [31:0] Prefetcher_io_out_bits_addr; // @[NutShell.scala 73:30]
  wire [2:0] Prefetcher_io_out_bits_size; // @[NutShell.scala 73:30]
  wire [3:0] Prefetcher_io_out_bits_cmd; // @[NutShell.scala 73:30]
  wire [7:0] Prefetcher_io_out_bits_wmask; // @[NutShell.scala 73:30]
  wire [63:0] Prefetcher_io_out_bits_wdata; // @[NutShell.scala 73:30]
  wire  Cache_clock; // @[Cache.scala 678:35]
  wire  Cache_reset; // @[Cache.scala 678:35]
  wire  Cache_io_in_req_ready; // @[Cache.scala 678:35]
  wire  Cache_io_in_req_valid; // @[Cache.scala 678:35]
  wire [31:0] Cache_io_in_req_bits_addr; // @[Cache.scala 678:35]
  wire [2:0] Cache_io_in_req_bits_size; // @[Cache.scala 678:35]
  wire [3:0] Cache_io_in_req_bits_cmd; // @[Cache.scala 678:35]
  wire [7:0] Cache_io_in_req_bits_wmask; // @[Cache.scala 678:35]
  wire [63:0] Cache_io_in_req_bits_wdata; // @[Cache.scala 678:35]
  wire  Cache_io_in_resp_valid; // @[Cache.scala 678:35]
  wire [3:0] Cache_io_in_resp_bits_cmd; // @[Cache.scala 678:35]
  wire [63:0] Cache_io_in_resp_bits_rdata; // @[Cache.scala 678:35]
  wire  Cache_io_out_mem_req_ready; // @[Cache.scala 678:35]
  wire  Cache_io_out_mem_req_valid; // @[Cache.scala 678:35]
  wire [31:0] Cache_io_out_mem_req_bits_addr; // @[Cache.scala 678:35]
  wire [3:0] Cache_io_out_mem_req_bits_cmd; // @[Cache.scala 678:35]
  wire [63:0] Cache_io_out_mem_req_bits_wdata; // @[Cache.scala 678:35]
  wire  Cache_io_out_mem_resp_valid; // @[Cache.scala 678:35]
  wire [3:0] Cache_io_out_mem_resp_bits_cmd; // @[Cache.scala 678:35]
  wire [63:0] Cache_io_out_mem_resp_bits_rdata; // @[Cache.scala 678:35]
  wire  memAddrMap_io_in_req_ready; // @[NutShell.scala 93:26]
  wire  memAddrMap_io_in_req_valid; // @[NutShell.scala 93:26]
  wire [31:0] memAddrMap_io_in_req_bits_addr; // @[NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_in_req_bits_cmd; // @[NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_in_req_bits_wdata; // @[NutShell.scala 93:26]
  wire  memAddrMap_io_in_resp_valid; // @[NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_in_resp_bits_cmd; // @[NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_in_resp_bits_rdata; // @[NutShell.scala 93:26]
  wire  memAddrMap_io_out_req_ready; // @[NutShell.scala 93:26]
  wire  memAddrMap_io_out_req_valid; // @[NutShell.scala 93:26]
  wire [31:0] memAddrMap_io_out_req_bits_addr; // @[NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_out_req_bits_cmd; // @[NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_out_req_bits_wdata; // @[NutShell.scala 93:26]
  wire  memAddrMap_io_out_resp_valid; // @[NutShell.scala 93:26]
  wire [3:0] memAddrMap_io_out_resp_bits_cmd; // @[NutShell.scala 93:26]
  wire [63:0] memAddrMap_io_out_resp_bits_rdata; // @[NutShell.scala 93:26]
  wire  SimpleBus2AXI4Converter_clock; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_reset; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_in_req_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_in_req_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_io_in_req_bits_addr; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_io_in_req_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_io_in_req_bits_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_in_resp_valid; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_io_in_resp_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_io_in_resp_bits_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_awready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_awvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_io_out_awaddr; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_io_out_awprot; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_awid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_awuser; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_io_out_awlen; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_io_out_awsize; // @[ToAXI4.scala 204:24]
  wire [1:0] SimpleBus2AXI4Converter_io_out_awburst; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_awlock; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_io_out_awcache; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_io_out_awqos; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_wready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_wvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_io_out_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_wlast; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_bvalid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_arready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_arvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_io_out_araddr; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_io_out_arprot; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_arid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_aruser; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_io_out_arlen; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_io_out_arsize; // @[ToAXI4.scala 204:24]
  wire [1:0] SimpleBus2AXI4Converter_io_out_arburst; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_arlock; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_io_out_arcache; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_io_out_arqos; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_rvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_io_out_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_io_out_rlast; // @[ToAXI4.scala 204:24]
  wire  mmioXbar_clock; // @[NutShell.scala 106:24]
  wire  mmioXbar_reset; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_in_req_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_in_req_valid; // @[NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_in_req_bits_addr; // @[NutShell.scala 106:24]
  wire [2:0] mmioXbar_io_in_req_bits_size; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_in_req_bits_cmd; // @[NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_in_req_bits_wmask; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_in_req_bits_wdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_in_resp_valid; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_in_resp_bits_cmd; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_in_resp_bits_rdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_req_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_req_valid; // @[NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_out_0_req_bits_addr; // @[NutShell.scala 106:24]
  wire [2:0] mmioXbar_io_out_0_req_bits_size; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_0_req_bits_cmd; // @[NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_out_0_req_bits_wmask; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_0_req_bits_wdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_resp_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_0_resp_valid; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_0_resp_bits_cmd; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_0_resp_bits_rdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_req_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_req_valid; // @[NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_out_1_req_bits_addr; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_1_req_bits_cmd; // @[NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_out_1_req_bits_wmask; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_1_req_bits_wdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_resp_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_1_resp_valid; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_1_resp_bits_rdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_req_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_req_valid; // @[NutShell.scala 106:24]
  wire [31:0] mmioXbar_io_out_2_req_bits_addr; // @[NutShell.scala 106:24]
  wire [3:0] mmioXbar_io_out_2_req_bits_cmd; // @[NutShell.scala 106:24]
  wire [7:0] mmioXbar_io_out_2_req_bits_wmask; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_2_req_bits_wdata; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_resp_ready; // @[NutShell.scala 106:24]
  wire  mmioXbar_io_out_2_resp_valid; // @[NutShell.scala 106:24]
  wire [63:0] mmioXbar_io_out_2_resp_bits_rdata; // @[NutShell.scala 106:24]
  wire  SimpleBus2AXI4Converter_1_clock; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_reset; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_in_req_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_in_req_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_1_io_in_req_bits_addr; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_1_io_in_req_bits_size; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_1_io_in_req_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_1_io_in_req_bits_wmask; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_1_io_in_req_bits_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_in_resp_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_in_resp_valid; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_1_io_in_resp_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_1_io_in_resp_bits_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_awready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_awvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_1_io_out_awaddr; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_1_io_out_awprot; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_awid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_awuser; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_1_io_out_awlen; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_1_io_out_awsize; // @[ToAXI4.scala 204:24]
  wire [1:0] SimpleBus2AXI4Converter_1_io_out_awburst; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_awlock; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_1_io_out_awcache; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_1_io_out_awqos; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_wready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_wvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_1_io_out_wdata; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_1_io_out_wstrb; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_wlast; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_bready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_bvalid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_arready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_arvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_1_io_out_araddr; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_1_io_out_arprot; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_arid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_aruser; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_1_io_out_arlen; // @[ToAXI4.scala 204:24]
  wire [2:0] SimpleBus2AXI4Converter_1_io_out_arsize; // @[ToAXI4.scala 204:24]
  wire [1:0] SimpleBus2AXI4Converter_1_io_out_arburst; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_arlock; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_1_io_out_arcache; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_1_io_out_arqos; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_rready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_rvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_1_io_out_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_1_io_out_rlast; // @[ToAXI4.scala 204:24]
  wire  clint_clock; // @[NutShell.scala 113:21]
  wire  clint_reset; // @[NutShell.scala 113:21]
  wire  clint_io__in_awready; // @[NutShell.scala 113:21]
  wire  clint_io__in_awvalid; // @[NutShell.scala 113:21]
  wire [31:0] clint_io__in_awaddr; // @[NutShell.scala 113:21]
  wire  clint_io__in_wready; // @[NutShell.scala 113:21]
  wire  clint_io__in_wvalid; // @[NutShell.scala 113:21]
  wire [63:0] clint_io__in_wdata; // @[NutShell.scala 113:21]
  wire [7:0] clint_io__in_wstrb; // @[NutShell.scala 113:21]
  wire  clint_io__in_bready; // @[NutShell.scala 113:21]
  wire  clint_io__in_bvalid; // @[NutShell.scala 113:21]
  wire  clint_io__in_arready; // @[NutShell.scala 113:21]
  wire  clint_io__in_arvalid; // @[NutShell.scala 113:21]
  wire [31:0] clint_io__in_araddr; // @[NutShell.scala 113:21]
  wire  clint_io__in_rready; // @[NutShell.scala 113:21]
  wire  clint_io__in_rvalid; // @[NutShell.scala 113:21]
  wire [63:0] clint_io__in_rdata; // @[NutShell.scala 113:21]
  wire  clint_io__extra_mtip; // @[NutShell.scala 113:21]
  wire  clint_io__extra_msip; // @[NutShell.scala 113:21]
  wire  clint_io_extra_mtip; // @[NutShell.scala 113:21]
  wire  clint_io_extra_msip; // @[NutShell.scala 113:21]
  wire  SimpleBus2AXI4Converter_2_clock; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_reset; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_in_req_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_in_req_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_2_io_in_req_bits_addr; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_2_io_in_req_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_2_io_in_req_bits_wmask; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_2_io_in_req_bits_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_in_resp_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_in_resp_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_2_io_in_resp_bits_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_awready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_awvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_2_io_out_awaddr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_wready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_wvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_2_io_out_wdata; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_2_io_out_wstrb; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_bready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_bvalid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_arready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_arvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_2_io_out_araddr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_rready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_2_io_out_rvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_2_io_out_rdata; // @[ToAXI4.scala 204:24]
  wire  plic_clock; // @[NutShell.scala 120:20]
  wire  plic_reset; // @[NutShell.scala 120:20]
  wire  plic_io__in_awready; // @[NutShell.scala 120:20]
  wire  plic_io__in_awvalid; // @[NutShell.scala 120:20]
  wire [31:0] plic_io__in_awaddr; // @[NutShell.scala 120:20]
  wire  plic_io__in_wready; // @[NutShell.scala 120:20]
  wire  plic_io__in_wvalid; // @[NutShell.scala 120:20]
  wire [63:0] plic_io__in_wdata; // @[NutShell.scala 120:20]
  wire [7:0] plic_io__in_wstrb; // @[NutShell.scala 120:20]
  wire  plic_io__in_bready; // @[NutShell.scala 120:20]
  wire  plic_io__in_bvalid; // @[NutShell.scala 120:20]
  wire  plic_io__in_arready; // @[NutShell.scala 120:20]
  wire  plic_io__in_arvalid; // @[NutShell.scala 120:20]
  wire [31:0] plic_io__in_araddr; // @[NutShell.scala 120:20]
  wire  plic_io__in_rready; // @[NutShell.scala 120:20]
  wire  plic_io__in_rvalid; // @[NutShell.scala 120:20]
  wire [63:0] plic_io__in_rdata; // @[NutShell.scala 120:20]
  wire [2:0] plic_io__extra_intrVec; // @[NutShell.scala 120:20]
  wire  plic_io__extra_meip_0; // @[NutShell.scala 120:20]
  wire  plic_io_extra_meip_0; // @[NutShell.scala 120:20]
  wire  SimpleBus2AXI4Converter_3_clock; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_reset; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_in_req_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_in_req_valid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_3_io_in_req_bits_addr; // @[ToAXI4.scala 204:24]
  wire [3:0] SimpleBus2AXI4Converter_3_io_in_req_bits_cmd; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_3_io_in_req_bits_wmask; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_3_io_in_req_bits_wdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_in_resp_ready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_in_resp_valid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_3_io_in_resp_bits_rdata; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_awready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_awvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_3_io_out_awaddr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_wready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_wvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_3_io_out_wdata; // @[ToAXI4.scala 204:24]
  wire [7:0] SimpleBus2AXI4Converter_3_io_out_wstrb; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_bready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_bvalid; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_arready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_arvalid; // @[ToAXI4.scala 204:24]
  wire [31:0] SimpleBus2AXI4Converter_3_io_out_araddr; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_rready; // @[ToAXI4.scala 204:24]
  wire  SimpleBus2AXI4Converter_3_io_out_rvalid; // @[ToAXI4.scala 204:24]
  wire [63:0] SimpleBus2AXI4Converter_3_io_out_rdata; // @[ToAXI4.scala 204:24]
  reg [2:0] _T_4; // @[NutShell.scala 122:47]
  reg [2:0] _T_5; // @[NutShell.scala 122:39]
  wire  ilaWBUvalid = nutcore_io_in_valid_0;
  wire  ilaWBUrfWen = nutcore_io_wb_rfWen;
  wire [4:0] ilaWBUrfDest = nutcore_io_wb_rfDest;
  wire [38:0] ilaWBUpc = nutcore_io_in_bits_decode_cf_pc;
  wire [63:0] _T_8 = {{25'd0}, ilaWBUpc};
  wire [63:0] _T_9 = {{63'd0}, ilaWBUvalid};
  wire [63:0] _T_10 = {{63'd0}, ilaWBUrfWen};
  wire [63:0] _T_11 = {{59'd0}, ilaWBUrfDest};
  NutCore nutcore ( // @[NutShell.scala 53:23]
    .clock(nutcore_clock),
    .reset(nutcore_reset),
    .io_imem_mem_req_ready(nutcore_io_imem_mem_req_ready),
    .io_imem_mem_req_valid(nutcore_io_imem_mem_req_valid),
    .io_imem_mem_req_bits_addr(nutcore_io_imem_mem_req_bits_addr),
    .io_imem_mem_req_bits_cmd(nutcore_io_imem_mem_req_bits_cmd),
    .io_imem_mem_req_bits_wdata(nutcore_io_imem_mem_req_bits_wdata),
    .io_imem_mem_resp_valid(nutcore_io_imem_mem_resp_valid),
    .io_imem_mem_resp_bits_cmd(nutcore_io_imem_mem_resp_bits_cmd),
    .io_imem_mem_resp_bits_rdata(nutcore_io_imem_mem_resp_bits_rdata),
    .io_dmem_mem_req_ready(nutcore_io_dmem_mem_req_ready),
    .io_dmem_mem_req_valid(nutcore_io_dmem_mem_req_valid),
    .io_dmem_mem_req_bits_addr(nutcore_io_dmem_mem_req_bits_addr),
    .io_dmem_mem_req_bits_cmd(nutcore_io_dmem_mem_req_bits_cmd),
    .io_dmem_mem_req_bits_wdata(nutcore_io_dmem_mem_req_bits_wdata),
    .io_dmem_mem_resp_valid(nutcore_io_dmem_mem_resp_valid),
    .io_dmem_mem_resp_bits_cmd(nutcore_io_dmem_mem_resp_bits_cmd),
    .io_dmem_mem_resp_bits_rdata(nutcore_io_dmem_mem_resp_bits_rdata),
    .io_dmem_coh_req_ready(nutcore_io_dmem_coh_req_ready),
    .io_dmem_coh_req_valid(nutcore_io_dmem_coh_req_valid),
    .io_dmem_coh_req_bits_addr(nutcore_io_dmem_coh_req_bits_addr),
    .io_dmem_coh_req_bits_wdata(nutcore_io_dmem_coh_req_bits_wdata),
    .io_dmem_coh_resp_valid(nutcore_io_dmem_coh_resp_valid),
    .io_dmem_coh_resp_bits_cmd(nutcore_io_dmem_coh_resp_bits_cmd),
    .io_dmem_coh_resp_bits_rdata(nutcore_io_dmem_coh_resp_bits_rdata),
    .io_mmio_req_ready(nutcore_io_mmio_req_ready),
    .io_mmio_req_valid(nutcore_io_mmio_req_valid),
    .io_mmio_req_bits_addr(nutcore_io_mmio_req_bits_addr),
    .io_mmio_req_bits_size(nutcore_io_mmio_req_bits_size),
    .io_mmio_req_bits_cmd(nutcore_io_mmio_req_bits_cmd),
    .io_mmio_req_bits_wmask(nutcore_io_mmio_req_bits_wmask),
    .io_mmio_req_bits_wdata(nutcore_io_mmio_req_bits_wdata),
    .io_mmio_resp_valid(nutcore_io_mmio_resp_valid),
    .io_mmio_resp_bits_cmd(nutcore_io_mmio_resp_bits_cmd),
    .io_mmio_resp_bits_rdata(nutcore_io_mmio_resp_bits_rdata),
    .io_frontend_req_ready(nutcore_io_frontend_req_ready),
    .io_frontend_req_valid(nutcore_io_frontend_req_valid),
    .io_frontend_req_bits_addr(nutcore_io_frontend_req_bits_addr),
    .io_frontend_req_bits_size(nutcore_io_frontend_req_bits_size),
    .io_frontend_req_bits_cmd(nutcore_io_frontend_req_bits_cmd),
    .io_frontend_req_bits_wmask(nutcore_io_frontend_req_bits_wmask),
    .io_frontend_req_bits_wdata(nutcore_io_frontend_req_bits_wdata),
    .io_frontend_resp_ready(nutcore_io_frontend_resp_ready),
    .io_frontend_resp_valid(nutcore_io_frontend_resp_valid),
    .io_frontend_resp_bits_cmd(nutcore_io_frontend_resp_bits_cmd),
    .io_frontend_resp_bits_rdata(nutcore_io_frontend_resp_bits_rdata),
    .perfCnts_2(nutcore_perfCnts_2),
    .io_in_bits_decode_cf_pc(nutcore_io_in_bits_decode_cf_pc),
    .io_wb_rfDest(nutcore_io_wb_rfDest),
    .io_extra_mtip(nutcore_io_extra_mtip),
    .io_extra_meip_0(nutcore_io_extra_meip_0),
    .io_wb_rfWen(nutcore_io_wb_rfWen),
    .io_wb_rfData(nutcore_io_wb_rfData),
    .io_extra_msip(nutcore_io_extra_msip),
    .io_in_valid_0(nutcore_io_in_valid_0)
  );
  CoherenceManager cohMg ( // @[NutShell.scala 54:21]
    .clock(cohMg_clock),
    .reset(cohMg_reset),
    .io_in_req_ready(cohMg_io_in_req_ready),
    .io_in_req_valid(cohMg_io_in_req_valid),
    .io_in_req_bits_addr(cohMg_io_in_req_bits_addr),
    .io_in_req_bits_cmd(cohMg_io_in_req_bits_cmd),
    .io_in_req_bits_wdata(cohMg_io_in_req_bits_wdata),
    .io_in_resp_valid(cohMg_io_in_resp_valid),
    .io_in_resp_bits_cmd(cohMg_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(cohMg_io_in_resp_bits_rdata),
    .io_out_mem_req_ready(cohMg_io_out_mem_req_ready),
    .io_out_mem_req_valid(cohMg_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(cohMg_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_cmd(cohMg_io_out_mem_req_bits_cmd),
    .io_out_mem_req_bits_wdata(cohMg_io_out_mem_req_bits_wdata),
    .io_out_mem_resp_ready(cohMg_io_out_mem_resp_ready),
    .io_out_mem_resp_valid(cohMg_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(cohMg_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(cohMg_io_out_mem_resp_bits_rdata),
    .io_out_coh_req_ready(cohMg_io_out_coh_req_ready),
    .io_out_coh_req_valid(cohMg_io_out_coh_req_valid),
    .io_out_coh_req_bits_addr(cohMg_io_out_coh_req_bits_addr),
    .io_out_coh_req_bits_wdata(cohMg_io_out_coh_req_bits_wdata),
    .io_out_coh_resp_ready(cohMg_io_out_coh_resp_ready),
    .io_out_coh_resp_valid(cohMg_io_out_coh_resp_valid),
    .io_out_coh_resp_bits_cmd(cohMg_io_out_coh_resp_bits_cmd),
    .io_out_coh_resp_bits_rdata(cohMg_io_out_coh_resp_bits_rdata)
  );
  SimpleBusCrossbarNto1 xbar ( // @[NutShell.scala 55:20]
    .clock(xbar_clock),
    .reset(xbar_reset),
    .io_in_0_req_ready(xbar_io_in_0_req_ready),
    .io_in_0_req_valid(xbar_io_in_0_req_valid),
    .io_in_0_req_bits_addr(xbar_io_in_0_req_bits_addr),
    .io_in_0_req_bits_cmd(xbar_io_in_0_req_bits_cmd),
    .io_in_0_req_bits_wmask(xbar_io_in_0_req_bits_wmask),
    .io_in_0_req_bits_wdata(xbar_io_in_0_req_bits_wdata),
    .io_in_0_resp_valid(xbar_io_in_0_resp_valid),
    .io_in_0_resp_bits_cmd(xbar_io_in_0_resp_bits_cmd),
    .io_in_0_resp_bits_rdata(xbar_io_in_0_resp_bits_rdata),
    .io_in_1_req_ready(xbar_io_in_1_req_ready),
    .io_in_1_req_valid(xbar_io_in_1_req_valid),
    .io_in_1_req_bits_addr(xbar_io_in_1_req_bits_addr),
    .io_in_1_req_bits_size(xbar_io_in_1_req_bits_size),
    .io_in_1_req_bits_cmd(xbar_io_in_1_req_bits_cmd),
    .io_in_1_req_bits_wmask(xbar_io_in_1_req_bits_wmask),
    .io_in_1_req_bits_wdata(xbar_io_in_1_req_bits_wdata),
    .io_in_1_resp_valid(xbar_io_in_1_resp_valid),
    .io_in_1_resp_bits_cmd(xbar_io_in_1_resp_bits_cmd),
    .io_in_1_resp_bits_rdata(xbar_io_in_1_resp_bits_rdata),
    .io_out_req_ready(xbar_io_out_req_ready),
    .io_out_req_valid(xbar_io_out_req_valid),
    .io_out_req_bits_addr(xbar_io_out_req_bits_addr),
    .io_out_req_bits_size(xbar_io_out_req_bits_size),
    .io_out_req_bits_cmd(xbar_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(xbar_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(xbar_io_out_req_bits_wdata),
    .io_out_resp_ready(xbar_io_out_resp_ready),
    .io_out_resp_valid(xbar_io_out_resp_valid),
    .io_out_resp_bits_cmd(xbar_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(xbar_io_out_resp_bits_rdata)
  );
  AXI42SimpleBusConverter axi2sb ( // @[NutShell.scala 61:22]
    .clock(axi2sb_clock),
    .reset(axi2sb_reset),
    .io_in_awready(axi2sb_io_in_awready),
    .io_in_awvalid(axi2sb_io_in_awvalid),
    .io_in_awaddr(axi2sb_io_in_awaddr),
    .io_in_awid(axi2sb_io_in_awid),
    .io_in_awlen(axi2sb_io_in_awlen),
    .io_in_awsize(axi2sb_io_in_awsize),
    .io_in_wready(axi2sb_io_in_wready),
    .io_in_wvalid(axi2sb_io_in_wvalid),
    .io_in_wdata(axi2sb_io_in_wdata),
    .io_in_wstrb(axi2sb_io_in_wstrb),
    .io_in_wlast(axi2sb_io_in_wlast),
    .io_in_bready(axi2sb_io_in_bready),
    .io_in_bvalid(axi2sb_io_in_bvalid),
    .io_in_arready(axi2sb_io_in_arready),
    .io_in_arvalid(axi2sb_io_in_arvalid),
    .io_in_araddr(axi2sb_io_in_araddr),
    .io_in_arid(axi2sb_io_in_arid),
    .io_in_arlen(axi2sb_io_in_arlen),
    .io_in_arsize(axi2sb_io_in_arsize),
    .io_in_rready(axi2sb_io_in_rready),
    .io_in_rvalid(axi2sb_io_in_rvalid),
    .io_in_rdata(axi2sb_io_in_rdata),
    .io_in_rlast(axi2sb_io_in_rlast),
    .io_in_rid(axi2sb_io_in_rid),
    .io_out_req_ready(axi2sb_io_out_req_ready),
    .io_out_req_valid(axi2sb_io_out_req_valid),
    .io_out_req_bits_addr(axi2sb_io_out_req_bits_addr),
    .io_out_req_bits_size(axi2sb_io_out_req_bits_size),
    .io_out_req_bits_cmd(axi2sb_io_out_req_bits_cmd),
    .io_out_req_bits_wmask(axi2sb_io_out_req_bits_wmask),
    .io_out_req_bits_wdata(axi2sb_io_out_req_bits_wdata),
    .io_out_resp_ready(axi2sb_io_out_resp_ready),
    .io_out_resp_valid(axi2sb_io_out_resp_valid),
    .io_out_resp_bits_cmd(axi2sb_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(axi2sb_io_out_resp_bits_rdata)
  );
  Prefetcher Prefetcher ( // @[NutShell.scala 73:30]
    .clock(Prefetcher_clock),
    .reset(Prefetcher_reset),
    .io_in_ready(Prefetcher_io_in_ready),
    .io_in_valid(Prefetcher_io_in_valid),
    .io_in_bits_addr(Prefetcher_io_in_bits_addr),
    .io_in_bits_size(Prefetcher_io_in_bits_size),
    .io_in_bits_cmd(Prefetcher_io_in_bits_cmd),
    .io_in_bits_wmask(Prefetcher_io_in_bits_wmask),
    .io_in_bits_wdata(Prefetcher_io_in_bits_wdata),
    .io_out_ready(Prefetcher_io_out_ready),
    .io_out_valid(Prefetcher_io_out_valid),
    .io_out_bits_addr(Prefetcher_io_out_bits_addr),
    .io_out_bits_size(Prefetcher_io_out_bits_size),
    .io_out_bits_cmd(Prefetcher_io_out_bits_cmd),
    .io_out_bits_wmask(Prefetcher_io_out_bits_wmask),
    .io_out_bits_wdata(Prefetcher_io_out_bits_wdata)
  );
  Cache_2 Cache ( // @[Cache.scala 678:35]
    .clock(Cache_clock),
    .reset(Cache_reset),
    .io_in_req_ready(Cache_io_in_req_ready),
    .io_in_req_valid(Cache_io_in_req_valid),
    .io_in_req_bits_addr(Cache_io_in_req_bits_addr),
    .io_in_req_bits_size(Cache_io_in_req_bits_size),
    .io_in_req_bits_cmd(Cache_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(Cache_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(Cache_io_in_req_bits_wdata),
    .io_in_resp_valid(Cache_io_in_resp_valid),
    .io_in_resp_bits_cmd(Cache_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(Cache_io_in_resp_bits_rdata),
    .io_out_mem_req_ready(Cache_io_out_mem_req_ready),
    .io_out_mem_req_valid(Cache_io_out_mem_req_valid),
    .io_out_mem_req_bits_addr(Cache_io_out_mem_req_bits_addr),
    .io_out_mem_req_bits_cmd(Cache_io_out_mem_req_bits_cmd),
    .io_out_mem_req_bits_wdata(Cache_io_out_mem_req_bits_wdata),
    .io_out_mem_resp_valid(Cache_io_out_mem_resp_valid),
    .io_out_mem_resp_bits_cmd(Cache_io_out_mem_resp_bits_cmd),
    .io_out_mem_resp_bits_rdata(Cache_io_out_mem_resp_bits_rdata)
  );
  SimpleBusAddressMapper memAddrMap ( // @[NutShell.scala 93:26]
    .io_in_req_ready(memAddrMap_io_in_req_ready),
    .io_in_req_valid(memAddrMap_io_in_req_valid),
    .io_in_req_bits_addr(memAddrMap_io_in_req_bits_addr),
    .io_in_req_bits_cmd(memAddrMap_io_in_req_bits_cmd),
    .io_in_req_bits_wdata(memAddrMap_io_in_req_bits_wdata),
    .io_in_resp_valid(memAddrMap_io_in_resp_valid),
    .io_in_resp_bits_cmd(memAddrMap_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(memAddrMap_io_in_resp_bits_rdata),
    .io_out_req_ready(memAddrMap_io_out_req_ready),
    .io_out_req_valid(memAddrMap_io_out_req_valid),
    .io_out_req_bits_addr(memAddrMap_io_out_req_bits_addr),
    .io_out_req_bits_cmd(memAddrMap_io_out_req_bits_cmd),
    .io_out_req_bits_wdata(memAddrMap_io_out_req_bits_wdata),
    .io_out_resp_valid(memAddrMap_io_out_resp_valid),
    .io_out_resp_bits_cmd(memAddrMap_io_out_resp_bits_cmd),
    .io_out_resp_bits_rdata(memAddrMap_io_out_resp_bits_rdata)
  );
  SimpleBus2AXI4Converter SimpleBus2AXI4Converter ( // @[ToAXI4.scala 204:24]
    .clock(SimpleBus2AXI4Converter_clock),
    .reset(SimpleBus2AXI4Converter_reset),
    .io_in_req_ready(SimpleBus2AXI4Converter_io_in_req_ready),
    .io_in_req_valid(SimpleBus2AXI4Converter_io_in_req_valid),
    .io_in_req_bits_addr(SimpleBus2AXI4Converter_io_in_req_bits_addr),
    .io_in_req_bits_cmd(SimpleBus2AXI4Converter_io_in_req_bits_cmd),
    .io_in_req_bits_wdata(SimpleBus2AXI4Converter_io_in_req_bits_wdata),
    .io_in_resp_valid(SimpleBus2AXI4Converter_io_in_resp_valid),
    .io_in_resp_bits_cmd(SimpleBus2AXI4Converter_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(SimpleBus2AXI4Converter_io_in_resp_bits_rdata),
    .io_out_awready(SimpleBus2AXI4Converter_io_out_awready),
    .io_out_awvalid(SimpleBus2AXI4Converter_io_out_awvalid),
    .io_out_awaddr(SimpleBus2AXI4Converter_io_out_awaddr),
    .io_out_awprot(SimpleBus2AXI4Converter_io_out_awprot),
    .io_out_awid(SimpleBus2AXI4Converter_io_out_awid),
    .io_out_awuser(SimpleBus2AXI4Converter_io_out_awuser),
    .io_out_awlen(SimpleBus2AXI4Converter_io_out_awlen),
    .io_out_awsize(SimpleBus2AXI4Converter_io_out_awsize),
    .io_out_awburst(SimpleBus2AXI4Converter_io_out_awburst),
    .io_out_awlock(SimpleBus2AXI4Converter_io_out_awlock),
    .io_out_awcache(SimpleBus2AXI4Converter_io_out_awcache),
    .io_out_awqos(SimpleBus2AXI4Converter_io_out_awqos),
    .io_out_wready(SimpleBus2AXI4Converter_io_out_wready),
    .io_out_wvalid(SimpleBus2AXI4Converter_io_out_wvalid),
    .io_out_wdata(SimpleBus2AXI4Converter_io_out_wdata),
    .io_out_wlast(SimpleBus2AXI4Converter_io_out_wlast),
    .io_out_bvalid(SimpleBus2AXI4Converter_io_out_bvalid),
    .io_out_arready(SimpleBus2AXI4Converter_io_out_arready),
    .io_out_arvalid(SimpleBus2AXI4Converter_io_out_arvalid),
    .io_out_araddr(SimpleBus2AXI4Converter_io_out_araddr),
    .io_out_arprot(SimpleBus2AXI4Converter_io_out_arprot),
    .io_out_arid(SimpleBus2AXI4Converter_io_out_arid),
    .io_out_aruser(SimpleBus2AXI4Converter_io_out_aruser),
    .io_out_arlen(SimpleBus2AXI4Converter_io_out_arlen),
    .io_out_arsize(SimpleBus2AXI4Converter_io_out_arsize),
    .io_out_arburst(SimpleBus2AXI4Converter_io_out_arburst),
    .io_out_arlock(SimpleBus2AXI4Converter_io_out_arlock),
    .io_out_arcache(SimpleBus2AXI4Converter_io_out_arcache),
    .io_out_arqos(SimpleBus2AXI4Converter_io_out_arqos),
    .io_out_rvalid(SimpleBus2AXI4Converter_io_out_rvalid),
    .io_out_rdata(SimpleBus2AXI4Converter_io_out_rdata),
    .io_out_rlast(SimpleBus2AXI4Converter_io_out_rlast)
  );
  SimpleBusCrossbar1toN mmioXbar ( // @[NutShell.scala 106:24]
    .clock(mmioXbar_clock),
    .reset(mmioXbar_reset),
    .io_in_req_ready(mmioXbar_io_in_req_ready),
    .io_in_req_valid(mmioXbar_io_in_req_valid),
    .io_in_req_bits_addr(mmioXbar_io_in_req_bits_addr),
    .io_in_req_bits_size(mmioXbar_io_in_req_bits_size),
    .io_in_req_bits_cmd(mmioXbar_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(mmioXbar_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(mmioXbar_io_in_req_bits_wdata),
    .io_in_resp_valid(mmioXbar_io_in_resp_valid),
    .io_in_resp_bits_cmd(mmioXbar_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(mmioXbar_io_in_resp_bits_rdata),
    .io_out_0_req_ready(mmioXbar_io_out_0_req_ready),
    .io_out_0_req_valid(mmioXbar_io_out_0_req_valid),
    .io_out_0_req_bits_addr(mmioXbar_io_out_0_req_bits_addr),
    .io_out_0_req_bits_size(mmioXbar_io_out_0_req_bits_size),
    .io_out_0_req_bits_cmd(mmioXbar_io_out_0_req_bits_cmd),
    .io_out_0_req_bits_wmask(mmioXbar_io_out_0_req_bits_wmask),
    .io_out_0_req_bits_wdata(mmioXbar_io_out_0_req_bits_wdata),
    .io_out_0_resp_ready(mmioXbar_io_out_0_resp_ready),
    .io_out_0_resp_valid(mmioXbar_io_out_0_resp_valid),
    .io_out_0_resp_bits_cmd(mmioXbar_io_out_0_resp_bits_cmd),
    .io_out_0_resp_bits_rdata(mmioXbar_io_out_0_resp_bits_rdata),
    .io_out_1_req_ready(mmioXbar_io_out_1_req_ready),
    .io_out_1_req_valid(mmioXbar_io_out_1_req_valid),
    .io_out_1_req_bits_addr(mmioXbar_io_out_1_req_bits_addr),
    .io_out_1_req_bits_cmd(mmioXbar_io_out_1_req_bits_cmd),
    .io_out_1_req_bits_wmask(mmioXbar_io_out_1_req_bits_wmask),
    .io_out_1_req_bits_wdata(mmioXbar_io_out_1_req_bits_wdata),
    .io_out_1_resp_ready(mmioXbar_io_out_1_resp_ready),
    .io_out_1_resp_valid(mmioXbar_io_out_1_resp_valid),
    .io_out_1_resp_bits_rdata(mmioXbar_io_out_1_resp_bits_rdata),
    .io_out_2_req_ready(mmioXbar_io_out_2_req_ready),
    .io_out_2_req_valid(mmioXbar_io_out_2_req_valid),
    .io_out_2_req_bits_addr(mmioXbar_io_out_2_req_bits_addr),
    .io_out_2_req_bits_cmd(mmioXbar_io_out_2_req_bits_cmd),
    .io_out_2_req_bits_wmask(mmioXbar_io_out_2_req_bits_wmask),
    .io_out_2_req_bits_wdata(mmioXbar_io_out_2_req_bits_wdata),
    .io_out_2_resp_ready(mmioXbar_io_out_2_resp_ready),
    .io_out_2_resp_valid(mmioXbar_io_out_2_resp_valid),
    .io_out_2_resp_bits_rdata(mmioXbar_io_out_2_resp_bits_rdata)
  );
  SimpleBus2AXI4Converter_1 SimpleBus2AXI4Converter_1 ( // @[ToAXI4.scala 204:24]
    .clock(SimpleBus2AXI4Converter_1_clock),
    .reset(SimpleBus2AXI4Converter_1_reset),
    .io_in_req_ready(SimpleBus2AXI4Converter_1_io_in_req_ready),
    .io_in_req_valid(SimpleBus2AXI4Converter_1_io_in_req_valid),
    .io_in_req_bits_addr(SimpleBus2AXI4Converter_1_io_in_req_bits_addr),
    .io_in_req_bits_size(SimpleBus2AXI4Converter_1_io_in_req_bits_size),
    .io_in_req_bits_cmd(SimpleBus2AXI4Converter_1_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(SimpleBus2AXI4Converter_1_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(SimpleBus2AXI4Converter_1_io_in_req_bits_wdata),
    .io_in_resp_ready(SimpleBus2AXI4Converter_1_io_in_resp_ready),
    .io_in_resp_valid(SimpleBus2AXI4Converter_1_io_in_resp_valid),
    .io_in_resp_bits_cmd(SimpleBus2AXI4Converter_1_io_in_resp_bits_cmd),
    .io_in_resp_bits_rdata(SimpleBus2AXI4Converter_1_io_in_resp_bits_rdata),
    .io_out_awready(SimpleBus2AXI4Converter_1_io_out_awready),
    .io_out_awvalid(SimpleBus2AXI4Converter_1_io_out_awvalid),
    .io_out_awaddr(SimpleBus2AXI4Converter_1_io_out_awaddr),
    .io_out_awprot(SimpleBus2AXI4Converter_1_io_out_awprot),
    .io_out_awid(SimpleBus2AXI4Converter_1_io_out_awid),
    .io_out_awuser(SimpleBus2AXI4Converter_1_io_out_awuser),
    .io_out_awlen(SimpleBus2AXI4Converter_1_io_out_awlen),
    .io_out_awsize(SimpleBus2AXI4Converter_1_io_out_awsize),
    .io_out_awburst(SimpleBus2AXI4Converter_1_io_out_awburst),
    .io_out_awlock(SimpleBus2AXI4Converter_1_io_out_awlock),
    .io_out_awcache(SimpleBus2AXI4Converter_1_io_out_awcache),
    .io_out_awqos(SimpleBus2AXI4Converter_1_io_out_awqos),
    .io_out_wready(SimpleBus2AXI4Converter_1_io_out_wready),
    .io_out_wvalid(SimpleBus2AXI4Converter_1_io_out_wvalid),
    .io_out_wdata(SimpleBus2AXI4Converter_1_io_out_wdata),
    .io_out_wstrb(SimpleBus2AXI4Converter_1_io_out_wstrb),
    .io_out_wlast(SimpleBus2AXI4Converter_1_io_out_wlast),
    .io_out_bready(SimpleBus2AXI4Converter_1_io_out_bready),
    .io_out_bvalid(SimpleBus2AXI4Converter_1_io_out_bvalid),
    .io_out_arready(SimpleBus2AXI4Converter_1_io_out_arready),
    .io_out_arvalid(SimpleBus2AXI4Converter_1_io_out_arvalid),
    .io_out_araddr(SimpleBus2AXI4Converter_1_io_out_araddr),
    .io_out_arprot(SimpleBus2AXI4Converter_1_io_out_arprot),
    .io_out_arid(SimpleBus2AXI4Converter_1_io_out_arid),
    .io_out_aruser(SimpleBus2AXI4Converter_1_io_out_aruser),
    .io_out_arlen(SimpleBus2AXI4Converter_1_io_out_arlen),
    .io_out_arsize(SimpleBus2AXI4Converter_1_io_out_arsize),
    .io_out_arburst(SimpleBus2AXI4Converter_1_io_out_arburst),
    .io_out_arlock(SimpleBus2AXI4Converter_1_io_out_arlock),
    .io_out_arcache(SimpleBus2AXI4Converter_1_io_out_arcache),
    .io_out_arqos(SimpleBus2AXI4Converter_1_io_out_arqos),
    .io_out_rready(SimpleBus2AXI4Converter_1_io_out_rready),
    .io_out_rvalid(SimpleBus2AXI4Converter_1_io_out_rvalid),
    .io_out_rdata(SimpleBus2AXI4Converter_1_io_out_rdata),
    .io_out_rlast(SimpleBus2AXI4Converter_1_io_out_rlast)
  );
  AXI4CLINT clint ( // @[NutShell.scala 113:21]
    .clock(clint_clock),
    .reset(clint_reset),
    .io__in_awready(clint_io__in_awready),
    .io__in_awvalid(clint_io__in_awvalid),
    .io__in_awaddr(clint_io__in_awaddr),
    .io__in_wready(clint_io__in_wready),
    .io__in_wvalid(clint_io__in_wvalid),
    .io__in_wdata(clint_io__in_wdata),
    .io__in_wstrb(clint_io__in_wstrb),
    .io__in_bready(clint_io__in_bready),
    .io__in_bvalid(clint_io__in_bvalid),
    .io__in_arready(clint_io__in_arready),
    .io__in_arvalid(clint_io__in_arvalid),
    .io__in_araddr(clint_io__in_araddr),
    .io__in_rready(clint_io__in_rready),
    .io__in_rvalid(clint_io__in_rvalid),
    .io__in_rdata(clint_io__in_rdata),
    .io__extra_mtip(clint_io__extra_mtip),
    .io__extra_msip(clint_io__extra_msip),
    .io_extra_mtip(clint_io_extra_mtip),
    .io_extra_msip(clint_io_extra_msip)
  );
  SimpleBus2AXI4Converter_2 SimpleBus2AXI4Converter_2 ( // @[ToAXI4.scala 204:24]
    .clock(SimpleBus2AXI4Converter_2_clock),
    .reset(SimpleBus2AXI4Converter_2_reset),
    .io_in_req_ready(SimpleBus2AXI4Converter_2_io_in_req_ready),
    .io_in_req_valid(SimpleBus2AXI4Converter_2_io_in_req_valid),
    .io_in_req_bits_addr(SimpleBus2AXI4Converter_2_io_in_req_bits_addr),
    .io_in_req_bits_cmd(SimpleBus2AXI4Converter_2_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(SimpleBus2AXI4Converter_2_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(SimpleBus2AXI4Converter_2_io_in_req_bits_wdata),
    .io_in_resp_ready(SimpleBus2AXI4Converter_2_io_in_resp_ready),
    .io_in_resp_valid(SimpleBus2AXI4Converter_2_io_in_resp_valid),
    .io_in_resp_bits_rdata(SimpleBus2AXI4Converter_2_io_in_resp_bits_rdata),
    .io_out_awready(SimpleBus2AXI4Converter_2_io_out_awready),
    .io_out_awvalid(SimpleBus2AXI4Converter_2_io_out_awvalid),
    .io_out_awaddr(SimpleBus2AXI4Converter_2_io_out_awaddr),
    .io_out_wready(SimpleBus2AXI4Converter_2_io_out_wready),
    .io_out_wvalid(SimpleBus2AXI4Converter_2_io_out_wvalid),
    .io_out_wdata(SimpleBus2AXI4Converter_2_io_out_wdata),
    .io_out_wstrb(SimpleBus2AXI4Converter_2_io_out_wstrb),
    .io_out_bready(SimpleBus2AXI4Converter_2_io_out_bready),
    .io_out_bvalid(SimpleBus2AXI4Converter_2_io_out_bvalid),
    .io_out_arready(SimpleBus2AXI4Converter_2_io_out_arready),
    .io_out_arvalid(SimpleBus2AXI4Converter_2_io_out_arvalid),
    .io_out_araddr(SimpleBus2AXI4Converter_2_io_out_araddr),
    .io_out_rready(SimpleBus2AXI4Converter_2_io_out_rready),
    .io_out_rvalid(SimpleBus2AXI4Converter_2_io_out_rvalid),
    .io_out_rdata(SimpleBus2AXI4Converter_2_io_out_rdata)
  );
  AXI4PLIC plic ( // @[NutShell.scala 120:20]
    .clock(plic_clock),
    .reset(plic_reset),
    .io__in_awready(plic_io__in_awready),
    .io__in_awvalid(plic_io__in_awvalid),
    .io__in_awaddr(plic_io__in_awaddr),
    .io__in_wready(plic_io__in_wready),
    .io__in_wvalid(plic_io__in_wvalid),
    .io__in_wdata(plic_io__in_wdata),
    .io__in_wstrb(plic_io__in_wstrb),
    .io__in_bready(plic_io__in_bready),
    .io__in_bvalid(plic_io__in_bvalid),
    .io__in_arready(plic_io__in_arready),
    .io__in_arvalid(plic_io__in_arvalid),
    .io__in_araddr(plic_io__in_araddr),
    .io__in_rready(plic_io__in_rready),
    .io__in_rvalid(plic_io__in_rvalid),
    .io__in_rdata(plic_io__in_rdata),
    .io__extra_intrVec(plic_io__extra_intrVec),
    .io__extra_meip_0(plic_io__extra_meip_0),
    .io_extra_meip_0(plic_io_extra_meip_0)
  );
  SimpleBus2AXI4Converter_2 SimpleBus2AXI4Converter_3 ( // @[ToAXI4.scala 204:24]
    .clock(SimpleBus2AXI4Converter_3_clock),
    .reset(SimpleBus2AXI4Converter_3_reset),
    .io_in_req_ready(SimpleBus2AXI4Converter_3_io_in_req_ready),
    .io_in_req_valid(SimpleBus2AXI4Converter_3_io_in_req_valid),
    .io_in_req_bits_addr(SimpleBus2AXI4Converter_3_io_in_req_bits_addr),
    .io_in_req_bits_cmd(SimpleBus2AXI4Converter_3_io_in_req_bits_cmd),
    .io_in_req_bits_wmask(SimpleBus2AXI4Converter_3_io_in_req_bits_wmask),
    .io_in_req_bits_wdata(SimpleBus2AXI4Converter_3_io_in_req_bits_wdata),
    .io_in_resp_ready(SimpleBus2AXI4Converter_3_io_in_resp_ready),
    .io_in_resp_valid(SimpleBus2AXI4Converter_3_io_in_resp_valid),
    .io_in_resp_bits_rdata(SimpleBus2AXI4Converter_3_io_in_resp_bits_rdata),
    .io_out_awready(SimpleBus2AXI4Converter_3_io_out_awready),
    .io_out_awvalid(SimpleBus2AXI4Converter_3_io_out_awvalid),
    .io_out_awaddr(SimpleBus2AXI4Converter_3_io_out_awaddr),
    .io_out_wready(SimpleBus2AXI4Converter_3_io_out_wready),
    .io_out_wvalid(SimpleBus2AXI4Converter_3_io_out_wvalid),
    .io_out_wdata(SimpleBus2AXI4Converter_3_io_out_wdata),
    .io_out_wstrb(SimpleBus2AXI4Converter_3_io_out_wstrb),
    .io_out_bready(SimpleBus2AXI4Converter_3_io_out_bready),
    .io_out_bvalid(SimpleBus2AXI4Converter_3_io_out_bvalid),
    .io_out_arready(SimpleBus2AXI4Converter_3_io_out_arready),
    .io_out_arvalid(SimpleBus2AXI4Converter_3_io_out_arvalid),
    .io_out_araddr(SimpleBus2AXI4Converter_3_io_out_araddr),
    .io_out_rready(SimpleBus2AXI4Converter_3_io_out_rready),
    .io_out_rvalid(SimpleBus2AXI4Converter_3_io_out_rvalid),
    .io_out_rdata(SimpleBus2AXI4Converter_3_io_out_rdata)
  );
  assign io_mem_awvalid = SimpleBus2AXI4Converter_io_out_awvalid; // @[NutShell.scala 95:10]
  assign io_mem_awaddr = SimpleBus2AXI4Converter_io_out_awaddr; // @[NutShell.scala 95:10]
  assign io_mem_awprot = SimpleBus2AXI4Converter_io_out_awprot; // @[NutShell.scala 95:10]
  assign io_mem_awid = SimpleBus2AXI4Converter_io_out_awid; // @[NutShell.scala 95:10]
  assign io_mem_awuser = SimpleBus2AXI4Converter_io_out_awuser; // @[NutShell.scala 95:10]
  assign io_mem_awlen = SimpleBus2AXI4Converter_io_out_awlen; // @[NutShell.scala 95:10]
  assign io_mem_awsize = SimpleBus2AXI4Converter_io_out_awsize; // @[NutShell.scala 95:10]
  assign io_mem_awburst = SimpleBus2AXI4Converter_io_out_awburst; // @[NutShell.scala 95:10]
  assign io_mem_awlock = SimpleBus2AXI4Converter_io_out_awlock; // @[NutShell.scala 95:10]
  assign io_mem_awcache = SimpleBus2AXI4Converter_io_out_awcache; // @[NutShell.scala 95:10]
  assign io_mem_awqos = SimpleBus2AXI4Converter_io_out_awqos; // @[NutShell.scala 95:10]
  assign io_mem_wvalid = SimpleBus2AXI4Converter_io_out_wvalid; // @[NutShell.scala 95:10]
  assign io_mem_wdata = SimpleBus2AXI4Converter_io_out_wdata; // @[NutShell.scala 95:10]
  assign io_mem_wstrb = 8'hff; // @[NutShell.scala 95:10]
  assign io_mem_wlast = SimpleBus2AXI4Converter_io_out_wlast; // @[NutShell.scala 95:10]
  assign io_mem_bready = 1'h1; // @[NutShell.scala 95:10]
  assign io_mem_arvalid = SimpleBus2AXI4Converter_io_out_arvalid; // @[NutShell.scala 95:10]
  assign io_mem_araddr = SimpleBus2AXI4Converter_io_out_araddr; // @[NutShell.scala 95:10]
  assign io_mem_arprot = 3'h1; // @[NutShell.scala 95:10]
  assign io_mem_arid = 1'h0; // @[NutShell.scala 95:10]
  assign io_mem_aruser = 1'h0; // @[NutShell.scala 95:10]
  assign io_mem_arlen = SimpleBus2AXI4Converter_io_out_arlen; // @[NutShell.scala 95:10]
  assign io_mem_arsize = 3'h3; // @[NutShell.scala 95:10]
  assign io_mem_arburst = 2'h2; // @[NutShell.scala 95:10]
  assign io_mem_arlock = 1'h0; // @[NutShell.scala 95:10]
  assign io_mem_arcache = 4'h0; // @[NutShell.scala 95:10]
  assign io_mem_arqos = 4'h0; // @[NutShell.scala 95:10]
  assign io_mem_rready = 1'h1; // @[NutShell.scala 95:10]
  assign io_mmio_awvalid = SimpleBus2AXI4Converter_1_io_out_awvalid; // @[NutShell.scala 110:33]
  assign io_mmio_awaddr = SimpleBus2AXI4Converter_1_io_out_awaddr; // @[NutShell.scala 110:33]
  assign io_mmio_awprot = SimpleBus2AXI4Converter_1_io_out_awprot; // @[NutShell.scala 110:33]
  assign io_mmio_awid = SimpleBus2AXI4Converter_1_io_out_awid; // @[NutShell.scala 110:33]
  assign io_mmio_awuser = SimpleBus2AXI4Converter_1_io_out_awuser; // @[NutShell.scala 110:33]
  assign io_mmio_awlen = SimpleBus2AXI4Converter_1_io_out_awlen; // @[NutShell.scala 110:33]
  assign io_mmio_awsize = SimpleBus2AXI4Converter_1_io_out_awsize; // @[NutShell.scala 110:33]
  assign io_mmio_awburst = SimpleBus2AXI4Converter_1_io_out_awburst; // @[NutShell.scala 110:33]
  assign io_mmio_awlock = SimpleBus2AXI4Converter_1_io_out_awlock; // @[NutShell.scala 110:33]
  assign io_mmio_awcache = SimpleBus2AXI4Converter_1_io_out_awcache; // @[NutShell.scala 110:33]
  assign io_mmio_awqos = SimpleBus2AXI4Converter_1_io_out_awqos; // @[NutShell.scala 110:33]
  assign io_mmio_wvalid = SimpleBus2AXI4Converter_1_io_out_wvalid; // @[NutShell.scala 110:33]
  assign io_mmio_wdata = SimpleBus2AXI4Converter_1_io_out_wdata; // @[NutShell.scala 110:33]
  assign io_mmio_wstrb = SimpleBus2AXI4Converter_1_io_out_wstrb; // @[NutShell.scala 110:33]
  assign io_mmio_wlast = SimpleBus2AXI4Converter_1_io_out_wlast; // @[NutShell.scala 110:33]
  assign io_mmio_bready = SimpleBus2AXI4Converter_1_io_out_bready; // @[NutShell.scala 110:33]
  assign io_mmio_arvalid = SimpleBus2AXI4Converter_1_io_out_arvalid; // @[NutShell.scala 110:33]
  assign io_mmio_araddr = SimpleBus2AXI4Converter_1_io_out_araddr; // @[NutShell.scala 110:33]
  assign io_mmio_arprot = 3'h1; // @[NutShell.scala 110:33]
  assign io_mmio_arid = 1'h0; // @[NutShell.scala 110:33]
  assign io_mmio_aruser = 1'h0; // @[NutShell.scala 110:33]
  assign io_mmio_arlen = SimpleBus2AXI4Converter_1_io_out_arlen; // @[NutShell.scala 110:33]
  assign io_mmio_arsize = SimpleBus2AXI4Converter_1_io_out_arsize; // @[NutShell.scala 110:33]
  assign io_mmio_arburst = 2'h1; // @[NutShell.scala 110:33]
  assign io_mmio_arlock = 1'h0; // @[NutShell.scala 110:33]
  assign io_mmio_arcache = 4'h0; // @[NutShell.scala 110:33]
  assign io_mmio_arqos = 4'h0; // @[NutShell.scala 110:33]
  assign io_mmio_rready = SimpleBus2AXI4Converter_1_io_out_rready; // @[NutShell.scala 110:33]
  assign io_frontend_awready = axi2sb_io_in_awready; // @[NutShell.scala 62:16]
  assign io_frontend_wready = axi2sb_io_in_wready; // @[NutShell.scala 62:16]
  assign io_frontend_bvalid = axi2sb_io_in_bvalid; // @[NutShell.scala 62:16]
  assign io_frontend_bresp = 2'h0; // @[NutShell.scala 62:16]
  assign io_frontend_bid = 1'h0; // @[NutShell.scala 62:16]
  assign io_frontend_buser = 1'h0; // @[NutShell.scala 62:16]
  assign io_frontend_arready = axi2sb_io_in_arready; // @[NutShell.scala 62:16]
  assign io_frontend_rvalid = axi2sb_io_in_rvalid; // @[NutShell.scala 62:16]
  assign io_frontend_rresp = 2'h0; // @[NutShell.scala 62:16]
  assign io_frontend_rdata = axi2sb_io_in_rdata; // @[NutShell.scala 62:16]
  assign io_frontend_rlast = axi2sb_io_in_rlast; // @[NutShell.scala 62:16]
  assign io_frontend_rid = axi2sb_io_in_rid[0]; // @[NutShell.scala 62:16]
  assign io_frontend_ruser = 1'h0; // @[NutShell.scala 62:16]
  assign io_ila_WBUpc = _T_8[38:0]; // @[NutShell.scala 132:12]
  assign io_ila_WBUvalid = _T_9[0]; // @[NutShell.scala 132:12]
  assign io_ila_WBUrfWen = _T_10[0]; // @[NutShell.scala 132:12]
  assign io_ila_WBUrfDest = _T_11[4:0]; // @[NutShell.scala 132:12]
  assign io_ila_WBUrfData = nutcore_io_wb_rfData; // @[NutShell.scala 132:12]
  assign io_ila_InstrCnt = nutcore_perfCnts_2; // @[NutShell.scala 132:12]
  assign nutcore_clock = clock;
  assign nutcore_reset = reset;
  assign nutcore_io_imem_mem_req_ready = cohMg_io_in_req_ready; // @[NutShell.scala 56:15]
  assign nutcore_io_imem_mem_resp_valid = cohMg_io_in_resp_valid; // @[NutShell.scala 56:15]
  assign nutcore_io_imem_mem_resp_bits_cmd = cohMg_io_in_resp_bits_cmd; // @[NutShell.scala 56:15]
  assign nutcore_io_imem_mem_resp_bits_rdata = cohMg_io_in_resp_bits_rdata; // @[NutShell.scala 56:15]
  assign nutcore_io_dmem_mem_req_ready = xbar_io_in_1_req_ready; // @[NutShell.scala 59:17]
  assign nutcore_io_dmem_mem_resp_valid = xbar_io_in_1_resp_valid; // @[NutShell.scala 59:17]
  assign nutcore_io_dmem_mem_resp_bits_cmd = xbar_io_in_1_resp_bits_cmd; // @[NutShell.scala 59:17]
  assign nutcore_io_dmem_mem_resp_bits_rdata = xbar_io_in_1_resp_bits_rdata; // @[NutShell.scala 59:17]
  assign nutcore_io_dmem_coh_req_valid = cohMg_io_out_coh_req_valid; // @[NutShell.scala 57:23]
  assign nutcore_io_dmem_coh_req_bits_addr = cohMg_io_out_coh_req_bits_addr; // @[NutShell.scala 57:23]
  assign nutcore_io_dmem_coh_req_bits_wdata = cohMg_io_out_coh_req_bits_wdata; // @[NutShell.scala 57:23]
  assign nutcore_io_mmio_req_ready = mmioXbar_io_in_req_ready; // @[NutShell.scala 107:18]
  assign nutcore_io_mmio_resp_valid = mmioXbar_io_in_resp_valid; // @[NutShell.scala 107:18]
  assign nutcore_io_mmio_resp_bits_cmd = mmioXbar_io_in_resp_bits_cmd; // @[NutShell.scala 107:18]
  assign nutcore_io_mmio_resp_bits_rdata = mmioXbar_io_in_resp_bits_rdata; // @[NutShell.scala 107:18]
  assign nutcore_io_frontend_req_valid = axi2sb_io_out_req_valid; // @[NutShell.scala 63:23]
  assign nutcore_io_frontend_req_bits_addr = axi2sb_io_out_req_bits_addr; // @[NutShell.scala 63:23]
  assign nutcore_io_frontend_req_bits_size = axi2sb_io_out_req_bits_size; // @[NutShell.scala 63:23]
  assign nutcore_io_frontend_req_bits_cmd = axi2sb_io_out_req_bits_cmd; // @[NutShell.scala 63:23]
  assign nutcore_io_frontend_req_bits_wmask = axi2sb_io_out_req_bits_wmask; // @[NutShell.scala 63:23]
  assign nutcore_io_frontend_req_bits_wdata = axi2sb_io_out_req_bits_wdata; // @[NutShell.scala 63:23]
  assign nutcore_io_frontend_resp_ready = axi2sb_io_out_resp_ready; // @[NutShell.scala 63:23]
  assign nutcore_io_extra_mtip = clint_io_extra_mtip;
  assign nutcore_io_extra_meip_0 = plic_io_extra_meip_0;
  assign nutcore_io_extra_msip = clint_io_extra_msip;
  assign cohMg_clock = clock;
  assign cohMg_reset = reset;
  assign cohMg_io_in_req_valid = nutcore_io_imem_mem_req_valid; // @[NutShell.scala 56:15]
  assign cohMg_io_in_req_bits_addr = nutcore_io_imem_mem_req_bits_addr; // @[NutShell.scala 56:15]
  assign cohMg_io_in_req_bits_cmd = nutcore_io_imem_mem_req_bits_cmd; // @[NutShell.scala 56:15]
  assign cohMg_io_in_req_bits_wdata = nutcore_io_imem_mem_req_bits_wdata; // @[NutShell.scala 56:15]
  assign cohMg_io_out_mem_req_ready = xbar_io_in_0_req_ready; // @[NutShell.scala 58:17]
  assign cohMg_io_out_mem_resp_valid = xbar_io_in_0_resp_valid; // @[NutShell.scala 58:17]
  assign cohMg_io_out_mem_resp_bits_cmd = xbar_io_in_0_resp_bits_cmd; // @[NutShell.scala 58:17]
  assign cohMg_io_out_mem_resp_bits_rdata = xbar_io_in_0_resp_bits_rdata; // @[NutShell.scala 58:17]
  assign cohMg_io_out_coh_req_ready = nutcore_io_dmem_coh_req_ready; // @[NutShell.scala 57:23]
  assign cohMg_io_out_coh_resp_valid = nutcore_io_dmem_coh_resp_valid; // @[NutShell.scala 57:23]
  assign cohMg_io_out_coh_resp_bits_cmd = nutcore_io_dmem_coh_resp_bits_cmd; // @[NutShell.scala 57:23]
  assign cohMg_io_out_coh_resp_bits_rdata = nutcore_io_dmem_coh_resp_bits_rdata; // @[NutShell.scala 57:23]
  assign xbar_clock = clock;
  assign xbar_reset = reset;
  assign xbar_io_in_0_req_valid = cohMg_io_out_mem_req_valid; // @[NutShell.scala 58:17]
  assign xbar_io_in_0_req_bits_addr = cohMg_io_out_mem_req_bits_addr; // @[NutShell.scala 58:17]
  assign xbar_io_in_0_req_bits_cmd = cohMg_io_out_mem_req_bits_cmd; // @[NutShell.scala 58:17]
  assign xbar_io_in_0_req_bits_wmask = 8'hff; // @[NutShell.scala 58:17]
  assign xbar_io_in_0_req_bits_wdata = cohMg_io_out_mem_req_bits_wdata; // @[NutShell.scala 58:17]
  assign xbar_io_in_1_req_valid = nutcore_io_dmem_mem_req_valid; // @[NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_addr = nutcore_io_dmem_mem_req_bits_addr; // @[NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_size = 3'h3; // @[NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_cmd = nutcore_io_dmem_mem_req_bits_cmd; // @[NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_wmask = 8'hff; // @[NutShell.scala 59:17]
  assign xbar_io_in_1_req_bits_wdata = nutcore_io_dmem_mem_req_bits_wdata; // @[NutShell.scala 59:17]
  assign xbar_io_out_req_ready = Prefetcher_io_in_ready; // @[ToMemPort.scala 51:18 NutShell.scala 75:24]
  assign xbar_io_out_resp_valid = Cache_io_in_resp_valid; // @[ToMemPort.scala 51:18 NutShell.scala 77:24]
  assign xbar_io_out_resp_bits_cmd = Cache_io_in_resp_bits_cmd; // @[ToMemPort.scala 51:18 NutShell.scala 77:24]
  assign xbar_io_out_resp_bits_rdata = Cache_io_in_resp_bits_rdata; // @[ToMemPort.scala 51:18 NutShell.scala 77:24]
  assign axi2sb_clock = clock;
  assign axi2sb_reset = reset;
  assign axi2sb_io_in_awvalid = io_frontend_awvalid; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_awaddr = io_frontend_awaddr; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_awid = {{17'd0}, io_frontend_awid}; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_awlen = io_frontend_awlen; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_awsize = io_frontend_awsize; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_wvalid = io_frontend_wvalid; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_wdata = io_frontend_wdata; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_wstrb = io_frontend_wstrb; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_wlast = io_frontend_wlast; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_bready = io_frontend_bready; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_arvalid = io_frontend_arvalid; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_araddr = io_frontend_araddr; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_arid = {{17'd0}, io_frontend_arid}; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_arlen = io_frontend_arlen; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_arsize = io_frontend_arsize; // @[NutShell.scala 62:16]
  assign axi2sb_io_in_rready = io_frontend_rready; // @[NutShell.scala 62:16]
  assign axi2sb_io_out_req_ready = nutcore_io_frontend_req_ready; // @[NutShell.scala 63:23]
  assign axi2sb_io_out_resp_valid = nutcore_io_frontend_resp_valid; // @[NutShell.scala 63:23]
  assign axi2sb_io_out_resp_bits_cmd = nutcore_io_frontend_resp_bits_cmd; // @[NutShell.scala 63:23]
  assign axi2sb_io_out_resp_bits_rdata = nutcore_io_frontend_resp_bits_rdata; // @[NutShell.scala 63:23]
  assign Prefetcher_clock = clock;
  assign Prefetcher_reset = reset;
  assign Prefetcher_io_in_valid = xbar_io_out_req_valid; // @[NutShell.scala 75:24]
  assign Prefetcher_io_in_bits_addr = xbar_io_out_req_bits_addr; // @[NutShell.scala 75:24]
  assign Prefetcher_io_in_bits_size = xbar_io_out_req_bits_size; // @[NutShell.scala 75:24]
  assign Prefetcher_io_in_bits_cmd = xbar_io_out_req_bits_cmd; // @[NutShell.scala 75:24]
  assign Prefetcher_io_in_bits_wmask = xbar_io_out_req_bits_wmask; // @[NutShell.scala 75:24]
  assign Prefetcher_io_in_bits_wdata = xbar_io_out_req_bits_wdata; // @[NutShell.scala 75:24]
  assign Prefetcher_io_out_ready = Cache_io_in_req_ready; // @[NutShell.scala 76:21]
  assign Cache_clock = clock;
  assign Cache_reset = reset;
  assign Cache_io_in_req_valid = Prefetcher_io_out_valid; // @[Cache.scala 684:17]
  assign Cache_io_in_req_bits_addr = Prefetcher_io_out_bits_addr; // @[Cache.scala 684:17]
  assign Cache_io_in_req_bits_size = Prefetcher_io_out_bits_size; // @[Cache.scala 684:17]
  assign Cache_io_in_req_bits_cmd = Prefetcher_io_out_bits_cmd; // @[Cache.scala 684:17]
  assign Cache_io_in_req_bits_wmask = Prefetcher_io_out_bits_wmask; // @[Cache.scala 684:17]
  assign Cache_io_in_req_bits_wdata = Prefetcher_io_out_bits_wdata; // @[Cache.scala 684:17]
  assign Cache_io_out_mem_req_ready = memAddrMap_io_in_req_ready; // @[NutShell.scala 81:16]
  assign Cache_io_out_mem_resp_valid = memAddrMap_io_in_resp_valid; // @[NutShell.scala 81:16]
  assign Cache_io_out_mem_resp_bits_cmd = memAddrMap_io_in_resp_bits_cmd; // @[NutShell.scala 81:16]
  assign Cache_io_out_mem_resp_bits_rdata = memAddrMap_io_in_resp_bits_rdata; // @[NutShell.scala 81:16]
  assign memAddrMap_io_in_req_valid = Cache_io_out_mem_req_valid; // @[NutShell.scala 94:20]
  assign memAddrMap_io_in_req_bits_addr = Cache_io_out_mem_req_bits_addr; // @[NutShell.scala 94:20]
  assign memAddrMap_io_in_req_bits_cmd = Cache_io_out_mem_req_bits_cmd; // @[NutShell.scala 94:20]
  assign memAddrMap_io_in_req_bits_wdata = Cache_io_out_mem_req_bits_wdata; // @[NutShell.scala 94:20]
  assign memAddrMap_io_out_req_ready = SimpleBus2AXI4Converter_io_in_req_ready; // @[ToAXI4.scala 205:18]
  assign memAddrMap_io_out_resp_valid = SimpleBus2AXI4Converter_io_in_resp_valid; // @[ToAXI4.scala 205:18]
  assign memAddrMap_io_out_resp_bits_cmd = SimpleBus2AXI4Converter_io_in_resp_bits_cmd; // @[ToAXI4.scala 205:18]
  assign memAddrMap_io_out_resp_bits_rdata = SimpleBus2AXI4Converter_io_in_resp_bits_rdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_clock = clock;
  assign SimpleBus2AXI4Converter_reset = reset;
  assign SimpleBus2AXI4Converter_io_in_req_valid = memAddrMap_io_out_req_valid; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_in_req_bits_addr = memAddrMap_io_out_req_bits_addr; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_in_req_bits_cmd = memAddrMap_io_out_req_bits_cmd; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_in_req_bits_wdata = memAddrMap_io_out_req_bits_wdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_io_out_awready = io_mem_awready; // @[NutShell.scala 95:10]
  assign SimpleBus2AXI4Converter_io_out_wready = io_mem_wready; // @[NutShell.scala 95:10]
  assign SimpleBus2AXI4Converter_io_out_bvalid = io_mem_bvalid; // @[NutShell.scala 95:10]
  assign SimpleBus2AXI4Converter_io_out_arready = io_mem_arready; // @[NutShell.scala 95:10]
  assign SimpleBus2AXI4Converter_io_out_rvalid = io_mem_rvalid; // @[NutShell.scala 95:10]
  assign SimpleBus2AXI4Converter_io_out_rdata = io_mem_rdata; // @[NutShell.scala 95:10]
  assign SimpleBus2AXI4Converter_io_out_rlast = io_mem_rlast; // @[NutShell.scala 95:10]
  assign mmioXbar_clock = clock;
  assign mmioXbar_reset = reset;
  assign mmioXbar_io_in_req_valid = nutcore_io_mmio_req_valid; // @[NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_addr = nutcore_io_mmio_req_bits_addr; // @[NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_size = nutcore_io_mmio_req_bits_size; // @[NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_cmd = nutcore_io_mmio_req_bits_cmd; // @[NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_wmask = nutcore_io_mmio_req_bits_wmask; // @[NutShell.scala 107:18]
  assign mmioXbar_io_in_req_bits_wdata = nutcore_io_mmio_req_bits_wdata; // @[NutShell.scala 107:18]
  assign mmioXbar_io_out_0_req_ready = SimpleBus2AXI4Converter_1_io_in_req_ready; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_0_resp_valid = SimpleBus2AXI4Converter_1_io_in_resp_valid; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_0_resp_bits_cmd = SimpleBus2AXI4Converter_1_io_in_resp_bits_cmd; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_0_resp_bits_rdata = SimpleBus2AXI4Converter_1_io_in_resp_bits_rdata; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_1_req_ready = SimpleBus2AXI4Converter_2_io_in_req_ready; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_1_resp_valid = SimpleBus2AXI4Converter_2_io_in_resp_valid; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_1_resp_bits_rdata = SimpleBus2AXI4Converter_2_io_in_resp_bits_rdata; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_2_req_ready = SimpleBus2AXI4Converter_3_io_in_req_ready; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_2_resp_valid = SimpleBus2AXI4Converter_3_io_in_resp_valid; // @[ToAXI4.scala 205:18]
  assign mmioXbar_io_out_2_resp_bits_rdata = SimpleBus2AXI4Converter_3_io_in_resp_bits_rdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_clock = clock;
  assign SimpleBus2AXI4Converter_1_reset = reset;
  assign SimpleBus2AXI4Converter_1_io_in_req_valid = mmioXbar_io_out_0_req_valid; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_req_bits_addr = mmioXbar_io_out_0_req_bits_addr; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_req_bits_size = mmioXbar_io_out_0_req_bits_size; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_req_bits_cmd = mmioXbar_io_out_0_req_bits_cmd; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_req_bits_wmask = mmioXbar_io_out_0_req_bits_wmask; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_req_bits_wdata = mmioXbar_io_out_0_req_bits_wdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_in_resp_ready = mmioXbar_io_out_0_resp_ready; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_1_io_out_awready = io_mmio_awready; // @[NutShell.scala 110:33]
  assign SimpleBus2AXI4Converter_1_io_out_wready = io_mmio_wready; // @[NutShell.scala 110:33]
  assign SimpleBus2AXI4Converter_1_io_out_bvalid = io_mmio_bvalid; // @[NutShell.scala 110:33]
  assign SimpleBus2AXI4Converter_1_io_out_arready = io_mmio_arready; // @[NutShell.scala 110:33]
  assign SimpleBus2AXI4Converter_1_io_out_rvalid = io_mmio_rvalid; // @[NutShell.scala 110:33]
  assign SimpleBus2AXI4Converter_1_io_out_rdata = io_mmio_rdata; // @[NutShell.scala 110:33]
  assign SimpleBus2AXI4Converter_1_io_out_rlast = io_mmio_rlast; // @[NutShell.scala 110:33]
  assign clint_clock = clock;
  assign clint_reset = reset;
  assign clint_io__in_awvalid = SimpleBus2AXI4Converter_2_io_out_awvalid; // @[NutShell.scala 114:15]
  assign clint_io__in_awaddr = SimpleBus2AXI4Converter_2_io_out_awaddr; // @[NutShell.scala 114:15]
  assign clint_io__in_wvalid = SimpleBus2AXI4Converter_2_io_out_wvalid; // @[NutShell.scala 114:15]
  assign clint_io__in_wdata = SimpleBus2AXI4Converter_2_io_out_wdata; // @[NutShell.scala 114:15]
  assign clint_io__in_wstrb = SimpleBus2AXI4Converter_2_io_out_wstrb; // @[NutShell.scala 114:15]
  assign clint_io__in_bready = SimpleBus2AXI4Converter_2_io_out_bready; // @[NutShell.scala 114:15]
  assign clint_io__in_arvalid = SimpleBus2AXI4Converter_2_io_out_arvalid; // @[NutShell.scala 114:15]
  assign clint_io__in_araddr = SimpleBus2AXI4Converter_2_io_out_araddr; // @[NutShell.scala 114:15]
  assign clint_io__in_rready = SimpleBus2AXI4Converter_2_io_out_rready; // @[NutShell.scala 114:15]
  assign SimpleBus2AXI4Converter_2_clock = clock;
  assign SimpleBus2AXI4Converter_2_reset = reset;
  assign SimpleBus2AXI4Converter_2_io_in_req_valid = mmioXbar_io_out_1_req_valid; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_req_bits_addr = mmioXbar_io_out_1_req_bits_addr; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_req_bits_cmd = mmioXbar_io_out_1_req_bits_cmd; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_req_bits_wmask = mmioXbar_io_out_1_req_bits_wmask; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_req_bits_wdata = mmioXbar_io_out_1_req_bits_wdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_in_resp_ready = mmioXbar_io_out_1_resp_ready; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_2_io_out_awready = clint_io__in_awready; // @[NutShell.scala 114:15]
  assign SimpleBus2AXI4Converter_2_io_out_wready = clint_io__in_wready; // @[NutShell.scala 114:15]
  assign SimpleBus2AXI4Converter_2_io_out_bvalid = clint_io__in_bvalid; // @[NutShell.scala 114:15]
  assign SimpleBus2AXI4Converter_2_io_out_arready = clint_io__in_arready; // @[NutShell.scala 114:15]
  assign SimpleBus2AXI4Converter_2_io_out_rvalid = clint_io__in_rvalid; // @[NutShell.scala 114:15]
  assign SimpleBus2AXI4Converter_2_io_out_rdata = clint_io__in_rdata; // @[NutShell.scala 114:15]
  assign plic_clock = clock;
  assign plic_reset = reset;
  assign plic_io__in_awvalid = SimpleBus2AXI4Converter_3_io_out_awvalid; // @[NutShell.scala 121:14]
  assign plic_io__in_awaddr = SimpleBus2AXI4Converter_3_io_out_awaddr; // @[NutShell.scala 121:14]
  assign plic_io__in_wvalid = SimpleBus2AXI4Converter_3_io_out_wvalid; // @[NutShell.scala 121:14]
  assign plic_io__in_wdata = SimpleBus2AXI4Converter_3_io_out_wdata; // @[NutShell.scala 121:14]
  assign plic_io__in_wstrb = SimpleBus2AXI4Converter_3_io_out_wstrb; // @[NutShell.scala 121:14]
  assign plic_io__in_bready = SimpleBus2AXI4Converter_3_io_out_bready; // @[NutShell.scala 121:14]
  assign plic_io__in_arvalid = SimpleBus2AXI4Converter_3_io_out_arvalid; // @[NutShell.scala 121:14]
  assign plic_io__in_araddr = SimpleBus2AXI4Converter_3_io_out_araddr; // @[NutShell.scala 121:14]
  assign plic_io__in_rready = SimpleBus2AXI4Converter_3_io_out_rready; // @[NutShell.scala 121:14]
  assign plic_io__extra_intrVec = _T_5; // @[NutShell.scala 122:29]
  assign SimpleBus2AXI4Converter_3_clock = clock;
  assign SimpleBus2AXI4Converter_3_reset = reset;
  assign SimpleBus2AXI4Converter_3_io_in_req_valid = mmioXbar_io_out_2_req_valid; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_3_io_in_req_bits_addr = mmioXbar_io_out_2_req_bits_addr; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_3_io_in_req_bits_cmd = mmioXbar_io_out_2_req_bits_cmd; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_3_io_in_req_bits_wmask = mmioXbar_io_out_2_req_bits_wmask; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_3_io_in_req_bits_wdata = mmioXbar_io_out_2_req_bits_wdata; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_3_io_in_resp_ready = mmioXbar_io_out_2_resp_ready; // @[ToAXI4.scala 205:18]
  assign SimpleBus2AXI4Converter_3_io_out_awready = plic_io__in_awready; // @[NutShell.scala 121:14]
  assign SimpleBus2AXI4Converter_3_io_out_wready = plic_io__in_wready; // @[NutShell.scala 121:14]
  assign SimpleBus2AXI4Converter_3_io_out_bvalid = plic_io__in_bvalid; // @[NutShell.scala 121:14]
  assign SimpleBus2AXI4Converter_3_io_out_arready = plic_io__in_arready; // @[NutShell.scala 121:14]
  assign SimpleBus2AXI4Converter_3_io_out_rvalid = plic_io__in_rvalid; // @[NutShell.scala 121:14]
  assign SimpleBus2AXI4Converter_3_io_out_rdata = plic_io__in_rdata; // @[NutShell.scala 121:14]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_4 = _RAND_0[2:0];
  _RAND_1 = {1{`RANDOM}};
  _T_5 = _RAND_1[2:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    _T_4 <= io_meip;
    _T_5 <= _T_4;
  end
endmodule
module VGACtrl(
  input         clock,
  input         reset,
  output        io_in_awready,
  input         io_in_awvalid,
  output        io_in_wready,
  input         io_in_wvalid,
  input         io_in_bready,
  output        io_in_bvalid,
  output        io_in_arready,
  input         io_in_arvalid,
  input  [31:0] io_in_araddr,
  input         io_in_rready,
  output        io_in_rvalid,
  output [63:0] io_in_rdata
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
`endif // RANDOMIZE_REG_INIT
  wire  _T_30 = io_in_arready & io_in_arvalid; // @[Decoupled.scala 40:37]
  wire  _T_31 = io_in_rready & io_in_rvalid; // @[Decoupled.scala 40:37]
  reg  r_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_31 ? 1'h0 : r_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_1 = _T_30 | _GEN_0; // @[StopWatch.scala 27:20]
  wire  _T_33 = ~r_busy; // @[AXI4Slave.scala 71:32]
  reg  ren; // @[AXI4Slave.scala 73:17]
  wire  _T_42 = _T_30 | r_busy; // @[AXI4Slave.scala 74:52]
  wire  _T_43 = ren & _T_42; // @[AXI4Slave.scala 74:35]
  reg  _T_45; // @[StopWatch.scala 24:20]
  wire  _GEN_2 = _T_31 ? 1'h0 : _T_45; // @[StopWatch.scala 26:19]
  wire  _GEN_3 = _T_43 | _GEN_2; // @[StopWatch.scala 27:20]
  wire  _T_46 = io_in_awready & io_in_awvalid; // @[Decoupled.scala 40:37]
  wire  _T_47 = io_in_bready & io_in_bvalid; // @[Decoupled.scala 40:37]
  reg  w_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_4 = _T_47 ? 1'h0 : w_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_5 = _T_46 | _GEN_4; // @[StopWatch.scala 27:20]
  wire  _T_50 = io_in_wready & io_in_wvalid; // @[Decoupled.scala 40:37]
  reg  _T_53; // @[StopWatch.scala 24:20]
  wire  _GEN_6 = _T_47 ? 1'h0 : _T_53; // @[StopWatch.scala 26:19]
  wire  _GEN_7 = _T_50 | _GEN_6; // @[StopWatch.scala 27:20]
  wire  _T_88 = 4'h0 == io_in_araddr[3:0]; // @[LookupTree.scala 24:34]
  wire  _T_89 = 4'h4 == io_in_araddr[3:0]; // @[LookupTree.scala 24:34]
  wire [31:0] _T_90 = _T_88 ? 32'h190012c : 32'h0; // @[Mux.scala 27:72]
  wire  _T_91 = _T_89 & _T_46; // @[Mux.scala 27:72]
  wire [31:0] _GEN_8 = {{31'd0}, _T_91}; // @[Mux.scala 27:72]
  wire [31:0] _T_92 = _T_90 | _GEN_8; // @[Mux.scala 27:72]
  assign io_in_awready = ~w_busy; // @[AXI4Slave.scala 94:15]
  assign io_in_wready = io_in_awvalid | w_busy; // @[AXI4Slave.scala 95:15]
  assign io_in_bvalid = _T_53; // @[AXI4Slave.scala 97:14]
  assign io_in_arready = io_in_rready | _T_33; // @[AXI4Slave.scala 71:15]
  assign io_in_rvalid = _T_45; // @[AXI4Slave.scala 74:14]
  assign io_in_rdata = {{32'd0}, _T_92}; // @[RegMap.scala 30:11]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  r_busy = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  ren = _RAND_1[0:0];
  _RAND_2 = {1{`RANDOM}};
  _T_45 = _RAND_2[0:0];
  _RAND_3 = {1{`RANDOM}};
  w_busy = _RAND_3[0:0];
  _RAND_4 = {1{`RANDOM}};
  _T_53 = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      r_busy <= 1'h0;
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin
      ren <= 1'h0;
    end else begin
      ren <= _T_30;
    end
    if (reset) begin
      _T_45 <= 1'h0;
    end else begin
      _T_45 <= _GEN_3;
    end
    if (reset) begin
      w_busy <= 1'h0;
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin
      _T_53 <= 1'h0;
    end else begin
      _T_53 <= _GEN_7;
    end
  end
endmodule
module AXI4RAM(
  input         clock,
  input         reset,
  output        io_in_awready,
  input         io_in_awvalid,
  input  [31:0] io_in_awaddr,
  output        io_in_wready,
  input         io_in_wvalid,
  input  [63:0] io_in_wdata,
  input  [7:0]  io_in_wstrb,
  input         io_in_bready,
  output        io_in_bvalid,
  output        io_in_arready,
  input         io_in_arvalid,
  input  [31:0] io_in_araddr,
  input         io_in_rready,
  output        io_in_rvalid,
  output [63:0] io_in_rdata
);
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_5;
  reg [31:0] _RAND_7;
  reg [31:0] _RAND_9;
  reg [31:0] _RAND_11;
  reg [31:0] _RAND_13;
  reg [31:0] _RAND_15;
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_6;
  reg [31:0] _RAND_8;
  reg [31:0] _RAND_10;
  reg [31:0] _RAND_12;
  reg [31:0] _RAND_14;
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_16;
  reg [31:0] _RAND_17;
  reg [31:0] _RAND_18;
  reg [31:0] _RAND_19;
  reg [31:0] _RAND_20;
  reg [63:0] _RAND_21;
`endif // RANDOMIZE_REG_INIT
  reg [7:0] _T_62_0 [0:59999]; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_0__T_85_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_0__T_85_addr; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_0__T_82_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_0__T_82_addr; // @[AXI4RAM.scala 61:18]
  wire  _T_62_0__T_82_mask; // @[AXI4RAM.scala 61:18]
  wire  _T_62_0__T_82_en; // @[AXI4RAM.scala 61:18]
  reg [7:0] _T_62_1 [0:59999]; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_1__T_85_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_1__T_85_addr; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_1__T_82_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_1__T_82_addr; // @[AXI4RAM.scala 61:18]
  wire  _T_62_1__T_82_mask; // @[AXI4RAM.scala 61:18]
  wire  _T_62_1__T_82_en; // @[AXI4RAM.scala 61:18]
  reg [7:0] _T_62_2 [0:59999]; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_2__T_85_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_2__T_85_addr; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_2__T_82_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_2__T_82_addr; // @[AXI4RAM.scala 61:18]
  wire  _T_62_2__T_82_mask; // @[AXI4RAM.scala 61:18]
  wire  _T_62_2__T_82_en; // @[AXI4RAM.scala 61:18]
  reg [7:0] _T_62_3 [0:59999]; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_3__T_85_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_3__T_85_addr; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_3__T_82_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_3__T_82_addr; // @[AXI4RAM.scala 61:18]
  wire  _T_62_3__T_82_mask; // @[AXI4RAM.scala 61:18]
  wire  _T_62_3__T_82_en; // @[AXI4RAM.scala 61:18]
  reg [7:0] _T_62_4 [0:59999]; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_4__T_85_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_4__T_85_addr; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_4__T_82_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_4__T_82_addr; // @[AXI4RAM.scala 61:18]
  wire  _T_62_4__T_82_mask; // @[AXI4RAM.scala 61:18]
  wire  _T_62_4__T_82_en; // @[AXI4RAM.scala 61:18]
  reg [7:0] _T_62_5 [0:59999]; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_5__T_85_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_5__T_85_addr; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_5__T_82_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_5__T_82_addr; // @[AXI4RAM.scala 61:18]
  wire  _T_62_5__T_82_mask; // @[AXI4RAM.scala 61:18]
  wire  _T_62_5__T_82_en; // @[AXI4RAM.scala 61:18]
  reg [7:0] _T_62_6 [0:59999]; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_6__T_85_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_6__T_85_addr; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_6__T_82_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_6__T_82_addr; // @[AXI4RAM.scala 61:18]
  wire  _T_62_6__T_82_mask; // @[AXI4RAM.scala 61:18]
  wire  _T_62_6__T_82_en; // @[AXI4RAM.scala 61:18]
  reg [7:0] _T_62_7 [0:59999]; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_7__T_85_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_7__T_85_addr; // @[AXI4RAM.scala 61:18]
  wire [7:0] _T_62_7__T_82_data; // @[AXI4RAM.scala 61:18]
  wire [15:0] _T_62_7__T_82_addr; // @[AXI4RAM.scala 61:18]
  wire  _T_62_7__T_82_mask; // @[AXI4RAM.scala 61:18]
  wire  _T_62_7__T_82_en; // @[AXI4RAM.scala 61:18]
  wire  _T_30 = io_in_arready & io_in_arvalid; // @[Decoupled.scala 40:37]
  reg  r_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = io_in_rvalid ? 1'h0 : r_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_1 = _T_30 | _GEN_0; // @[StopWatch.scala 27:20]
  reg  ren; // @[AXI4Slave.scala 73:17]
  wire  _T_42 = _T_30 | r_busy; // @[AXI4Slave.scala 74:52]
  wire  _T_43 = ren & _T_42; // @[AXI4Slave.scala 74:35]
  reg  _T_45; // @[StopWatch.scala 24:20]
  wire  _GEN_2 = io_in_rvalid ? 1'h0 : _T_45; // @[StopWatch.scala 26:19]
  wire  _GEN_3 = _T_43 | _GEN_2; // @[StopWatch.scala 27:20]
  wire  _T_46 = io_in_awready & io_in_awvalid; // @[Decoupled.scala 40:37]
  wire  _T_47 = io_in_bready & io_in_bvalid; // @[Decoupled.scala 40:37]
  reg  w_busy; // @[StopWatch.scala 24:20]
  wire  _GEN_4 = _T_47 ? 1'h0 : w_busy; // @[StopWatch.scala 26:19]
  wire  _GEN_5 = _T_46 | _GEN_4; // @[StopWatch.scala 27:20]
  wire  _T_50 = io_in_wready & io_in_wvalid; // @[Decoupled.scala 40:37]
  reg  _T_53; // @[StopWatch.scala 24:20]
  wire  _GEN_6 = _T_47 ? 1'h0 : _T_53; // @[StopWatch.scala 26:19]
  wire  _GEN_7 = _T_50 | _GEN_6; // @[StopWatch.scala 27:20]
  wire [31:0] _T_54 = io_in_awaddr & 32'h7ffff; // @[AXI4RAM.scala 44:33]
  wire [29:0] _T_56 = {{1'd0}, _T_54[31:3]}; // @[AXI4RAM.scala 47:27]
  wire [28:0] wIdx = _T_56[28:0]; // @[AXI4RAM.scala 47:27]
  wire [31:0] _T_57 = io_in_araddr & 32'h7ffff; // @[AXI4RAM.scala 44:33]
  wire [29:0] _T_59 = {{1'd0}, _T_57[31:3]}; // @[AXI4RAM.scala 48:27]
  wire [28:0] rIdx = _T_59[28:0]; // @[AXI4RAM.scala 48:27]
  wire  _T_61 = wIdx < 29'hea60; // @[AXI4RAM.scala 45:32]
  wire [63:0] rdata = {_T_62_7__T_85_data,_T_62_6__T_85_data,_T_62_5__T_85_data,_T_62_4__T_85_data,_T_62_3__T_85_data,_T_62_2__T_85_data,_T_62_1__T_85_data,_T_62_0__T_85_data}; // @[Cat.scala 29:58]
  reg [63:0] _T_92; // @[Reg.scala 15:16]
  assign _T_62_0__T_85_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_0__T_85_data = _T_62_0[_T_62_0__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `else
  assign _T_62_0__T_85_data = _T_62_0__T_85_addr >= 16'hea60 ? _RAND_1[7:0] : _T_62_0[_T_62_0__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_0__T_82_data = io_in_wdata[7:0];
  assign _T_62_0__T_82_addr = wIdx[15:0];
  assign _T_62_0__T_82_mask = io_in_wstrb[0];
  assign _T_62_0__T_82_en = _T_50 & _T_61;
  assign _T_62_1__T_85_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_1__T_85_data = _T_62_1[_T_62_1__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `else
  assign _T_62_1__T_85_data = _T_62_1__T_85_addr >= 16'hea60 ? _RAND_3[7:0] : _T_62_1[_T_62_1__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_1__T_82_data = io_in_wdata[15:8];
  assign _T_62_1__T_82_addr = wIdx[15:0];
  assign _T_62_1__T_82_mask = io_in_wstrb[1];
  assign _T_62_1__T_82_en = _T_50 & _T_61;
  assign _T_62_2__T_85_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_2__T_85_data = _T_62_2[_T_62_2__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `else
  assign _T_62_2__T_85_data = _T_62_2__T_85_addr >= 16'hea60 ? _RAND_5[7:0] : _T_62_2[_T_62_2__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_2__T_82_data = io_in_wdata[23:16];
  assign _T_62_2__T_82_addr = wIdx[15:0];
  assign _T_62_2__T_82_mask = io_in_wstrb[2];
  assign _T_62_2__T_82_en = _T_50 & _T_61;
  assign _T_62_3__T_85_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_3__T_85_data = _T_62_3[_T_62_3__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `else
  assign _T_62_3__T_85_data = _T_62_3__T_85_addr >= 16'hea60 ? _RAND_7[7:0] : _T_62_3[_T_62_3__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_3__T_82_data = io_in_wdata[31:24];
  assign _T_62_3__T_82_addr = wIdx[15:0];
  assign _T_62_3__T_82_mask = io_in_wstrb[3];
  assign _T_62_3__T_82_en = _T_50 & _T_61;
  assign _T_62_4__T_85_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_4__T_85_data = _T_62_4[_T_62_4__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `else
  assign _T_62_4__T_85_data = _T_62_4__T_85_addr >= 16'hea60 ? _RAND_9[7:0] : _T_62_4[_T_62_4__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_4__T_82_data = io_in_wdata[39:32];
  assign _T_62_4__T_82_addr = wIdx[15:0];
  assign _T_62_4__T_82_mask = io_in_wstrb[4];
  assign _T_62_4__T_82_en = _T_50 & _T_61;
  assign _T_62_5__T_85_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_5__T_85_data = _T_62_5[_T_62_5__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `else
  assign _T_62_5__T_85_data = _T_62_5__T_85_addr >= 16'hea60 ? _RAND_11[7:0] : _T_62_5[_T_62_5__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_5__T_82_data = io_in_wdata[47:40];
  assign _T_62_5__T_82_addr = wIdx[15:0];
  assign _T_62_5__T_82_mask = io_in_wstrb[5];
  assign _T_62_5__T_82_en = _T_50 & _T_61;
  assign _T_62_6__T_85_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_6__T_85_data = _T_62_6[_T_62_6__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `else
  assign _T_62_6__T_85_data = _T_62_6__T_85_addr >= 16'hea60 ? _RAND_13[7:0] : _T_62_6[_T_62_6__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_6__T_82_data = io_in_wdata[55:48];
  assign _T_62_6__T_82_addr = wIdx[15:0];
  assign _T_62_6__T_82_mask = io_in_wstrb[6];
  assign _T_62_6__T_82_en = _T_50 & _T_61;
  assign _T_62_7__T_85_addr = rIdx[15:0];
  `ifndef RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_7__T_85_data = _T_62_7[_T_62_7__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `else
  assign _T_62_7__T_85_data = _T_62_7__T_85_addr >= 16'hea60 ? _RAND_15[7:0] : _T_62_7[_T_62_7__T_85_addr]; // @[AXI4RAM.scala 61:18]
  `endif // RANDOMIZE_GARBAGE_ASSIGN
  assign _T_62_7__T_82_data = io_in_wdata[63:56];
  assign _T_62_7__T_82_addr = wIdx[15:0];
  assign _T_62_7__T_82_mask = io_in_wstrb[7];
  assign _T_62_7__T_82_en = _T_50 & _T_61;
  assign io_in_awready = ~w_busy; // @[AXI4Slave.scala 94:15]
  assign io_in_wready = io_in_awvalid | w_busy; // @[AXI4Slave.scala 95:15]
  assign io_in_bvalid = _T_53; // @[AXI4Slave.scala 97:14]
  assign io_in_arready = 1'h1; // @[AXI4Slave.scala 71:15]
  assign io_in_rvalid = _T_45; // @[AXI4Slave.scala 74:14]
  assign io_in_rdata = _T_92; // @[AXI4RAM.scala 69:18]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_GARBAGE_ASSIGN
  _RAND_1 = {1{`RANDOM}};
  _RAND_3 = {1{`RANDOM}};
  _RAND_5 = {1{`RANDOM}};
  _RAND_7 = {1{`RANDOM}};
  _RAND_9 = {1{`RANDOM}};
  _RAND_11 = {1{`RANDOM}};
  _RAND_13 = {1{`RANDOM}};
  _RAND_15 = {1{`RANDOM}};
`endif // RANDOMIZE_GARBAGE_ASSIGN
`ifdef RANDOMIZE_MEM_INIT
  _RAND_0 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    _T_62_0[initvar] = _RAND_0[7:0];
  _RAND_2 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    _T_62_1[initvar] = _RAND_2[7:0];
  _RAND_4 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    _T_62_2[initvar] = _RAND_4[7:0];
  _RAND_6 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    _T_62_3[initvar] = _RAND_6[7:0];
  _RAND_8 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    _T_62_4[initvar] = _RAND_8[7:0];
  _RAND_10 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    _T_62_5[initvar] = _RAND_10[7:0];
  _RAND_12 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    _T_62_6[initvar] = _RAND_12[7:0];
  _RAND_14 = {1{`RANDOM}};
  for (initvar = 0; initvar < 60000; initvar = initvar+1)
    _T_62_7[initvar] = _RAND_14[7:0];
`endif // RANDOMIZE_MEM_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  r_busy = _RAND_16[0:0];
  _RAND_17 = {1{`RANDOM}};
  ren = _RAND_17[0:0];
  _RAND_18 = {1{`RANDOM}};
  _T_45 = _RAND_18[0:0];
  _RAND_19 = {1{`RANDOM}};
  w_busy = _RAND_19[0:0];
  _RAND_20 = {1{`RANDOM}};
  _T_53 = _RAND_20[0:0];
  _RAND_21 = {2{`RANDOM}};
  _T_92 = _RAND_21[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if(_T_62_0__T_82_en & _T_62_0__T_82_mask) begin
      _T_62_0[_T_62_0__T_82_addr] <= _T_62_0__T_82_data; // @[AXI4RAM.scala 61:18]
    end
    if(_T_62_1__T_82_en & _T_62_1__T_82_mask) begin
      _T_62_1[_T_62_1__T_82_addr] <= _T_62_1__T_82_data; // @[AXI4RAM.scala 61:18]
    end
    if(_T_62_2__T_82_en & _T_62_2__T_82_mask) begin
      _T_62_2[_T_62_2__T_82_addr] <= _T_62_2__T_82_data; // @[AXI4RAM.scala 61:18]
    end
    if(_T_62_3__T_82_en & _T_62_3__T_82_mask) begin
      _T_62_3[_T_62_3__T_82_addr] <= _T_62_3__T_82_data; // @[AXI4RAM.scala 61:18]
    end
    if(_T_62_4__T_82_en & _T_62_4__T_82_mask) begin
      _T_62_4[_T_62_4__T_82_addr] <= _T_62_4__T_82_data; // @[AXI4RAM.scala 61:18]
    end
    if(_T_62_5__T_82_en & _T_62_5__T_82_mask) begin
      _T_62_5[_T_62_5__T_82_addr] <= _T_62_5__T_82_data; // @[AXI4RAM.scala 61:18]
    end
    if(_T_62_6__T_82_en & _T_62_6__T_82_mask) begin
      _T_62_6[_T_62_6__T_82_addr] <= _T_62_6__T_82_data; // @[AXI4RAM.scala 61:18]
    end
    if(_T_62_7__T_82_en & _T_62_7__T_82_mask) begin
      _T_62_7[_T_62_7__T_82_addr] <= _T_62_7__T_82_data; // @[AXI4RAM.scala 61:18]
    end
    if (reset) begin
      r_busy <= 1'h0;
    end else begin
      r_busy <= _GEN_1;
    end
    if (reset) begin
      ren <= 1'h0;
    end else begin
      ren <= _T_30;
    end
    if (reset) begin
      _T_45 <= 1'h0;
    end else begin
      _T_45 <= _GEN_3;
    end
    if (reset) begin
      w_busy <= 1'h0;
    end else begin
      w_busy <= _GEN_5;
    end
    if (reset) begin
      _T_53 <= 1'h0;
    end else begin
      _T_53 <= _GEN_7;
    end
    if (ren) begin
      _T_92 <= rdata;
    end
  end
endmodule
module AXI4VGA(
  input         clock,
  input         reset,
  output        io_in_fb_awready,
  input         io_in_fb_awvalid,
  input  [31:0] io_in_fb_awaddr,
  input  [2:0]  io_in_fb_awprot,
  output        io_in_fb_wready,
  input         io_in_fb_wvalid,
  input  [63:0] io_in_fb_wdata,
  input  [7:0]  io_in_fb_wstrb,
  input         io_in_fb_bready,
  output        io_in_fb_bvalid,
  output [1:0]  io_in_fb_bresp,
  output        io_in_fb_arready,
  input         io_in_fb_arvalid,
  input  [31:0] io_in_fb_araddr,
  input  [2:0]  io_in_fb_arprot,
  input         io_in_fb_rready,
  output        io_in_fb_rvalid,
  output [1:0]  io_in_fb_rresp,
  output [63:0] io_in_fb_rdata,
  output        io_in_ctrl_awready,
  input         io_in_ctrl_awvalid,
  input  [31:0] io_in_ctrl_awaddr,
  input  [2:0]  io_in_ctrl_awprot,
  output        io_in_ctrl_wready,
  input         io_in_ctrl_wvalid,
  input  [63:0] io_in_ctrl_wdata,
  input  [7:0]  io_in_ctrl_wstrb,
  input         io_in_ctrl_bready,
  output        io_in_ctrl_bvalid,
  output [1:0]  io_in_ctrl_bresp,
  output        io_in_ctrl_arready,
  input         io_in_ctrl_arvalid,
  input  [31:0] io_in_ctrl_araddr,
  input  [2:0]  io_in_ctrl_arprot,
  input         io_in_ctrl_rready,
  output        io_in_ctrl_rvalid,
  output [1:0]  io_in_ctrl_rresp,
  output [63:0] io_in_ctrl_rdata,
  output [23:0] io_vga_rgb,
  output        io_vga_hsync,
  output        io_vga_vsync,
  output        io_vga_valid
);
`ifdef RANDOMIZE_REG_INIT
  reg [31:0] _RAND_0;
  reg [31:0] _RAND_1;
  reg [31:0] _RAND_2;
  reg [31:0] _RAND_3;
  reg [31:0] _RAND_4;
  reg [31:0] _RAND_5;
  reg [63:0] _RAND_6;
`endif // RANDOMIZE_REG_INIT
  wire  ctrl_clock; // @[AXI4VGA.scala 125:20]
  wire  ctrl_reset; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_awready; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_awvalid; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_wready; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_wvalid; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_bready; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_bvalid; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_arready; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_arvalid; // @[AXI4VGA.scala 125:20]
  wire [31:0] ctrl_io_in_araddr; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_rready; // @[AXI4VGA.scala 125:20]
  wire  ctrl_io_in_rvalid; // @[AXI4VGA.scala 125:20]
  wire [63:0] ctrl_io_in_rdata; // @[AXI4VGA.scala 125:20]
  wire  fb_clock; // @[AXI4VGA.scala 127:18]
  wire  fb_reset; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_awready; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_awvalid; // @[AXI4VGA.scala 127:18]
  wire [31:0] fb_io_in_awaddr; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_wready; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_wvalid; // @[AXI4VGA.scala 127:18]
  wire [63:0] fb_io_in_wdata; // @[AXI4VGA.scala 127:18]
  wire [7:0] fb_io_in_wstrb; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_bready; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_bvalid; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_arready; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_arvalid; // @[AXI4VGA.scala 127:18]
  wire [31:0] fb_io_in_araddr; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_rready; // @[AXI4VGA.scala 127:18]
  wire  fb_io_in_rvalid; // @[AXI4VGA.scala 127:18]
  wire [63:0] fb_io_in_rdata; // @[AXI4VGA.scala 127:18]
  wire  _T = io_in_fb_arready & io_in_fb_arvalid; // @[Decoupled.scala 40:37]
  wire  _T_1 = io_in_fb_rready & io_in_fb_rvalid; // @[Decoupled.scala 40:37]
  reg  _T_2; // @[StopWatch.scala 24:20]
  wire  _GEN_0 = _T_1 ? 1'h0 : _T_2; // @[StopWatch.scala 26:19]
  wire  _GEN_1 = _T | _GEN_0; // @[StopWatch.scala 27:20]
  reg [10:0] hCounter; // @[Counter.scala 29:33]
  wire  hFinish = hCounter == 11'h41f; // @[Counter.scala 38:24]
  wire [10:0] _T_5 = hCounter + 11'h1; // @[Counter.scala 39:22]
  reg [9:0] vCounter; // @[Counter.scala 29:33]
  wire  _T_6 = vCounter == 10'h273; // @[Counter.scala 38:24]
  wire [9:0] _T_8 = vCounter + 10'h1; // @[Counter.scala 39:22]
  wire  _T_11 = hCounter >= 11'ha8; // @[AXI4VGA.scala 138:51]
  wire  _T_12 = hCounter < 11'h3c8; // @[AXI4VGA.scala 138:69]
  wire  hInRange = _T_11 & _T_12; // @[AXI4VGA.scala 138:63]
  wire  _T_13 = vCounter >= 10'h5; // @[AXI4VGA.scala 138:51]
  wire  _T_14 = vCounter < 10'h25d; // @[AXI4VGA.scala 138:69]
  wire  vInRange = _T_13 & _T_14; // @[AXI4VGA.scala 138:63]
  wire  hCounterIsOdd = hCounter[0]; // @[AXI4VGA.scala 150:31]
  wire  hCounterIs2 = hCounter[1:0] == 2'h2; // @[AXI4VGA.scala 151:35]
  wire  vCounterIsOdd = vCounter[0]; // @[AXI4VGA.scala 152:31]
  wire  _T_17 = hCounter >= 11'ha7; // @[AXI4VGA.scala 138:51]
  wire  _T_18 = hCounter < 11'h3c7; // @[AXI4VGA.scala 138:69]
  wire  _T_19 = _T_17 & _T_18; // @[AXI4VGA.scala 138:63]
  wire  _T_20 = _T_19 & vInRange; // @[AXI4VGA.scala 155:66]
  wire  nextPixel = _T_20 & hCounterIsOdd; // @[AXI4VGA.scala 155:78]
  wire  _T_21 = ~vCounterIsOdd; // @[AXI4VGA.scala 156:44]
  wire  _T_22 = nextPixel & _T_21; // @[AXI4VGA.scala 156:41]
  reg [16:0] fbPixelAddrV0; // @[Counter.scala 29:33]
  wire  _T_24 = fbPixelAddrV0 == 17'h1d4bf; // @[Counter.scala 38:24]
  wire [16:0] _T_26 = fbPixelAddrV0 + 17'h1; // @[Counter.scala 39:22]
  wire  _T_27 = nextPixel & vCounterIsOdd; // @[AXI4VGA.scala 157:41]
  reg [16:0] fbPixelAddrV1; // @[Counter.scala 29:33]
  wire  _T_29 = fbPixelAddrV1 == 17'h1d4bf; // @[Counter.scala 38:24]
  wire [16:0] _T_31 = fbPixelAddrV1 + 17'h1; // @[Counter.scala 39:22]
  wire [16:0] _T_32 = vCounterIsOdd ? fbPixelAddrV1 : fbPixelAddrV0; // @[AXI4VGA.scala 161:35]
  wire [18:0] _T_33 = {_T_32,2'h0}; // @[Cat.scala 29:58]
  reg  _T_34; // @[AXI4VGA.scala 162:31]
  wire  _T_36 = fb_io_in_rready & fb_io_in_rvalid; // @[Decoupled.scala 40:37]
  reg [63:0] _T_38; // @[Reg.scala 27:20]
  wire [63:0] _GEN_14 = _T_36 ? fb_io_in_rdata : _T_38; // @[Reg.scala 28:19]
  wire [31:0] color = hCounter[1] ? _GEN_14[63:32] : _GEN_14[31:0]; // @[AXI4VGA.scala 167:23]
  VGACtrl ctrl ( // @[AXI4VGA.scala 125:20]
    .clock(ctrl_clock),
    .reset(ctrl_reset),
    .io_in_awready(ctrl_io_in_awready),
    .io_in_awvalid(ctrl_io_in_awvalid),
    .io_in_wready(ctrl_io_in_wready),
    .io_in_wvalid(ctrl_io_in_wvalid),
    .io_in_bready(ctrl_io_in_bready),
    .io_in_bvalid(ctrl_io_in_bvalid),
    .io_in_arready(ctrl_io_in_arready),
    .io_in_arvalid(ctrl_io_in_arvalid),
    .io_in_araddr(ctrl_io_in_araddr),
    .io_in_rready(ctrl_io_in_rready),
    .io_in_rvalid(ctrl_io_in_rvalid),
    .io_in_rdata(ctrl_io_in_rdata)
  );
  AXI4RAM fb ( // @[AXI4VGA.scala 127:18]
    .clock(fb_clock),
    .reset(fb_reset),
    .io_in_awready(fb_io_in_awready),
    .io_in_awvalid(fb_io_in_awvalid),
    .io_in_awaddr(fb_io_in_awaddr),
    .io_in_wready(fb_io_in_wready),
    .io_in_wvalid(fb_io_in_wvalid),
    .io_in_wdata(fb_io_in_wdata),
    .io_in_wstrb(fb_io_in_wstrb),
    .io_in_bready(fb_io_in_bready),
    .io_in_bvalid(fb_io_in_bvalid),
    .io_in_arready(fb_io_in_arready),
    .io_in_arvalid(fb_io_in_arvalid),
    .io_in_araddr(fb_io_in_araddr),
    .io_in_rready(fb_io_in_rready),
    .io_in_rvalid(fb_io_in_rvalid),
    .io_in_rdata(fb_io_in_rdata)
  );
  assign io_in_fb_awready = fb_io_in_awready; // @[AXI4VGA.scala 130:15]
  assign io_in_fb_wready = fb_io_in_wready; // @[AXI4VGA.scala 131:14]
  assign io_in_fb_bvalid = fb_io_in_bvalid; // @[AXI4VGA.scala 132:14]
  assign io_in_fb_bresp = 2'h0; // @[AXI4VGA.scala 132:14]
  assign io_in_fb_arready = 1'h1; // @[AXI4VGA.scala 133:21]
  assign io_in_fb_rvalid = _T_2; // @[AXI4VGA.scala 136:20]
  assign io_in_fb_rresp = 2'h0; // @[AXI4VGA.scala 135:24]
  assign io_in_fb_rdata = 64'h0; // @[AXI4VGA.scala 134:24]
  assign io_in_ctrl_awready = ctrl_io_in_awready; // @[AXI4VGA.scala 126:14]
  assign io_in_ctrl_wready = ctrl_io_in_wready; // @[AXI4VGA.scala 126:14]
  assign io_in_ctrl_bvalid = ctrl_io_in_bvalid; // @[AXI4VGA.scala 126:14]
  assign io_in_ctrl_bresp = 2'h0; // @[AXI4VGA.scala 126:14]
  assign io_in_ctrl_arready = ctrl_io_in_arready; // @[AXI4VGA.scala 126:14]
  assign io_in_ctrl_rvalid = ctrl_io_in_rvalid; // @[AXI4VGA.scala 126:14]
  assign io_in_ctrl_rresp = 2'h0; // @[AXI4VGA.scala 126:14]
  assign io_in_ctrl_rdata = ctrl_io_in_rdata; // @[AXI4VGA.scala 126:14]
  assign io_vga_rgb = io_vga_valid ? color[23:0] : 24'h0; // @[AXI4VGA.scala 168:14]
  assign io_vga_hsync = hCounter >= 11'h28; // @[AXI4VGA.scala 143:16]
  assign io_vga_vsync = vCounter >= 10'h1; // @[AXI4VGA.scala 144:16]
  assign io_vga_valid = hInRange & vInRange; // @[AXI4VGA.scala 148:16]
  assign ctrl_clock = clock;
  assign ctrl_reset = reset;
  assign ctrl_io_in_awvalid = io_in_ctrl_awvalid; // @[AXI4VGA.scala 126:14]
  assign ctrl_io_in_wvalid = io_in_ctrl_wvalid; // @[AXI4VGA.scala 126:14]
  assign ctrl_io_in_bready = io_in_ctrl_bready; // @[AXI4VGA.scala 126:14]
  assign ctrl_io_in_arvalid = io_in_ctrl_arvalid; // @[AXI4VGA.scala 126:14]
  assign ctrl_io_in_araddr = io_in_ctrl_araddr; // @[AXI4VGA.scala 126:14]
  assign ctrl_io_in_rready = io_in_ctrl_rready; // @[AXI4VGA.scala 126:14]
  assign fb_clock = clock;
  assign fb_reset = reset;
  assign fb_io_in_awvalid = io_in_fb_awvalid; // @[AXI4VGA.scala 130:15]
  assign fb_io_in_awaddr = io_in_fb_awaddr; // @[AXI4VGA.scala 130:15]
  assign fb_io_in_wvalid = io_in_fb_wvalid; // @[AXI4VGA.scala 131:14]
  assign fb_io_in_wdata = io_in_fb_wdata; // @[AXI4VGA.scala 131:14]
  assign fb_io_in_wstrb = io_in_fb_wstrb; // @[AXI4VGA.scala 131:14]
  assign fb_io_in_bready = io_in_fb_bready; // @[AXI4VGA.scala 132:14]
  assign fb_io_in_arvalid = _T_34 & hCounterIs2; // @[AXI4VGA.scala 162:21]
  assign fb_io_in_araddr = {{13'd0}, _T_33}; // @[AXI4VGA.scala 161:25]
  assign fb_io_in_rready = 1'h1; // @[AXI4VGA.scala 164:20]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE_MEM_INIT
  integer initvar;
`endif
`ifndef SYNTHESIS
`ifdef FIRRTL_BEFORE_INITIAL
`FIRRTL_BEFORE_INITIAL
`endif
initial begin
  `ifdef RANDOMIZE
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      `ifdef RANDOMIZE_DELAY
        #`RANDOMIZE_DELAY begin end
      `else
        #0.002 begin end
      `endif
    `endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  _T_2 = _RAND_0[0:0];
  _RAND_1 = {1{`RANDOM}};
  hCounter = _RAND_1[10:0];
  _RAND_2 = {1{`RANDOM}};
  vCounter = _RAND_2[9:0];
  _RAND_3 = {1{`RANDOM}};
  fbPixelAddrV0 = _RAND_3[16:0];
  _RAND_4 = {1{`RANDOM}};
  fbPixelAddrV1 = _RAND_4[16:0];
  _RAND_5 = {1{`RANDOM}};
  _T_34 = _RAND_5[0:0];
  _RAND_6 = {2{`RANDOM}};
  _T_38 = _RAND_6[63:0];
`endif // RANDOMIZE_REG_INIT
  `endif // RANDOMIZE
end // initial
`ifdef FIRRTL_AFTER_INITIAL
`FIRRTL_AFTER_INITIAL
`endif
`endif // SYNTHESIS
  always @(posedge clock) begin
    if (reset) begin
      _T_2 <= 1'h0;
    end else begin
      _T_2 <= _GEN_1;
    end
    if (reset) begin
      hCounter <= 11'h0;
    end else if (hFinish) begin
      hCounter <= 11'h0;
    end else begin
      hCounter <= _T_5;
    end
    if (reset) begin
      vCounter <= 10'h0;
    end else if (hFinish) begin
      if (_T_6) begin
        vCounter <= 10'h0;
      end else begin
        vCounter <= _T_8;
      end
    end
    if (reset) begin
      fbPixelAddrV0 <= 17'h0;
    end else if (_T_22) begin
      if (_T_24) begin
        fbPixelAddrV0 <= 17'h0;
      end else begin
        fbPixelAddrV0 <= _T_26;
      end
    end
    if (reset) begin
      fbPixelAddrV1 <= 17'h0;
    end else if (_T_27) begin
      if (_T_29) begin
        fbPixelAddrV1 <= 17'h0;
      end else begin
        fbPixelAddrV1 <= _T_31;
      end
    end
    _T_34 <= _T_20 & hCounterIsOdd;
    if (reset) begin
      _T_38 <= 64'h0;
    end else if (_T_36) begin
      _T_38 <= fb_io_in_rdata;
    end
  end
endmodule
module Top(
  input   clock,
  input   reset
);
  wire  nutshell_clock; // @[TopMain.scala 28:24]
  wire  nutshell_reset; // @[TopMain.scala 28:24]
  wire  nutshell_io_mem_awready; // @[TopMain.scala 28:24]
  wire  nutshell_io_mem_awvalid; // @[TopMain.scala 28:24]
  wire [31:0] nutshell_io_mem_awaddr; // @[TopMain.scala 28:24]
  wire [2:0] nutshell_io_mem_awprot; // @[TopMain.scala 28:24]
  wire  nutshell_io_mem_awid; // @[TopMain.scala 28:24]
  wire  nutshell_io_mem_awuser; // @[TopMain.scala 28:24]
  wire [7:0] nutshell_io_mem_awlen; // @[TopMain.scala 28:24]
  wire [2:0] nutshell_io_mem_awsize; // @[TopMain.scala 28:24]
  wire [1:0] nutshell_io_mem_awburst; // @[TopMain.scala 28:24]
  wire  nutshell_io_mem_awlock; // @[TopMain.scala 28:24]
  wire [3:0] nutshell_io_mem_awcache; // @[TopMain.scala 28:24]
  wire [3:0] nutshell_io_mem_awqos; // @[TopMain.scala 28:24]
  wire  nutshell_io_mem_wready; // @[TopMain.scala 28:24]
  wire  nutshell_io_mem_wvalid; // @[TopMain.scala 28:24]
  wire [63:0] nutshell_io_mem_wdata; // @[TopMain.scala 28:24]
  wire [7:0] nutshell_io_mem_wstrb; // @[TopMain.scala 28:24]
  wire  nutshell_io_mem_wlast; // @[TopMain.scala 28:24]
  wire  nutshell_io_mem_bready; // @[TopMain.scala 28:24]
  wire  nutshell_io_mem_bvalid; // @[TopMain.scala 28:24]
  wire [1:0] nutshell_io_mem_bresp; // @[TopMain.scala 28:24]
  wire  nutshell_io_mem_bid; // @[TopMain.scala 28:24]
  wire  nutshell_io_mem_buser; // @[TopMain.scala 28:24]
  wire  nutshell_io_mem_arready; // @[TopMain.scala 28:24]
  wire  nutshell_io_mem_arvalid; // @[TopMain.scala 28:24]
  wire [31:0] nutshell_io_mem_araddr; // @[TopMain.scala 28:24]
  wire [2:0] nutshell_io_mem_arprot; // @[TopMain.scala 28:24]
  wire  nutshell_io_mem_arid; // @[TopMain.scala 28:24]
  wire  nutshell_io_mem_aruser; // @[TopMain.scala 28:24]
  wire [7:0] nutshell_io_mem_arlen; // @[TopMain.scala 28:24]
  wire [2:0] nutshell_io_mem_arsize; // @[TopMain.scala 28:24]
  wire [1:0] nutshell_io_mem_arburst; // @[TopMain.scala 28:24]
  wire  nutshell_io_mem_arlock; // @[TopMain.scala 28:24]
  wire [3:0] nutshell_io_mem_arcache; // @[TopMain.scala 28:24]
  wire [3:0] nutshell_io_mem_arqos; // @[TopMain.scala 28:24]
  wire  nutshell_io_mem_rready; // @[TopMain.scala 28:24]
  wire  nutshell_io_mem_rvalid; // @[TopMain.scala 28:24]
  wire [1:0] nutshell_io_mem_rresp; // @[TopMain.scala 28:24]
  wire [63:0] nutshell_io_mem_rdata; // @[TopMain.scala 28:24]
  wire  nutshell_io_mem_rlast; // @[TopMain.scala 28:24]
  wire  nutshell_io_mem_rid; // @[TopMain.scala 28:24]
  wire  nutshell_io_mem_ruser; // @[TopMain.scala 28:24]
  wire  nutshell_io_mmio_awready; // @[TopMain.scala 28:24]
  wire  nutshell_io_mmio_awvalid; // @[TopMain.scala 28:24]
  wire [31:0] nutshell_io_mmio_awaddr; // @[TopMain.scala 28:24]
  wire [2:0] nutshell_io_mmio_awprot; // @[TopMain.scala 28:24]
  wire  nutshell_io_mmio_awid; // @[TopMain.scala 28:24]
  wire  nutshell_io_mmio_awuser; // @[TopMain.scala 28:24]
  wire [7:0] nutshell_io_mmio_awlen; // @[TopMain.scala 28:24]
  wire [2:0] nutshell_io_mmio_awsize; // @[TopMain.scala 28:24]
  wire [1:0] nutshell_io_mmio_awburst; // @[TopMain.scala 28:24]
  wire  nutshell_io_mmio_awlock; // @[TopMain.scala 28:24]
  wire [3:0] nutshell_io_mmio_awcache; // @[TopMain.scala 28:24]
  wire [3:0] nutshell_io_mmio_awqos; // @[TopMain.scala 28:24]
  wire  nutshell_io_mmio_wready; // @[TopMain.scala 28:24]
  wire  nutshell_io_mmio_wvalid; // @[TopMain.scala 28:24]
  wire [63:0] nutshell_io_mmio_wdata; // @[TopMain.scala 28:24]
  wire [7:0] nutshell_io_mmio_wstrb; // @[TopMain.scala 28:24]
  wire  nutshell_io_mmio_wlast; // @[TopMain.scala 28:24]
  wire  nutshell_io_mmio_bready; // @[TopMain.scala 28:24]
  wire  nutshell_io_mmio_bvalid; // @[TopMain.scala 28:24]
  wire [1:0] nutshell_io_mmio_bresp; // @[TopMain.scala 28:24]
  wire  nutshell_io_mmio_bid; // @[TopMain.scala 28:24]
  wire  nutshell_io_mmio_buser; // @[TopMain.scala 28:24]
  wire  nutshell_io_mmio_arready; // @[TopMain.scala 28:24]
  wire  nutshell_io_mmio_arvalid; // @[TopMain.scala 28:24]
  wire [31:0] nutshell_io_mmio_araddr; // @[TopMain.scala 28:24]
  wire [2:0] nutshell_io_mmio_arprot; // @[TopMain.scala 28:24]
  wire  nutshell_io_mmio_arid; // @[TopMain.scala 28:24]
  wire  nutshell_io_mmio_aruser; // @[TopMain.scala 28:24]
  wire [7:0] nutshell_io_mmio_arlen; // @[TopMain.scala 28:24]
  wire [2:0] nutshell_io_mmio_arsize; // @[TopMain.scala 28:24]
  wire [1:0] nutshell_io_mmio_arburst; // @[TopMain.scala 28:24]
  wire  nutshell_io_mmio_arlock; // @[TopMain.scala 28:24]
  wire [3:0] nutshell_io_mmio_arcache; // @[TopMain.scala 28:24]
  wire [3:0] nutshell_io_mmio_arqos; // @[TopMain.scala 28:24]
  wire  nutshell_io_mmio_rready; // @[TopMain.scala 28:24]
  wire  nutshell_io_mmio_rvalid; // @[TopMain.scala 28:24]
  wire [1:0] nutshell_io_mmio_rresp; // @[TopMain.scala 28:24]
  wire [63:0] nutshell_io_mmio_rdata; // @[TopMain.scala 28:24]
  wire  nutshell_io_mmio_rlast; // @[TopMain.scala 28:24]
  wire  nutshell_io_mmio_rid; // @[TopMain.scala 28:24]
  wire  nutshell_io_mmio_ruser; // @[TopMain.scala 28:24]
  wire  nutshell_io_frontend_awready; // @[TopMain.scala 28:24]
  wire  nutshell_io_frontend_awvalid; // @[TopMain.scala 28:24]
  wire [31:0] nutshell_io_frontend_awaddr; // @[TopMain.scala 28:24]
  wire [2:0] nutshell_io_frontend_awprot; // @[TopMain.scala 28:24]
  wire  nutshell_io_frontend_awid; // @[TopMain.scala 28:24]
  wire  nutshell_io_frontend_awuser; // @[TopMain.scala 28:24]
  wire [7:0] nutshell_io_frontend_awlen; // @[TopMain.scala 28:24]
  wire [2:0] nutshell_io_frontend_awsize; // @[TopMain.scala 28:24]
  wire [1:0] nutshell_io_frontend_awburst; // @[TopMain.scala 28:24]
  wire  nutshell_io_frontend_awlock; // @[TopMain.scala 28:24]
  wire [3:0] nutshell_io_frontend_awcache; // @[TopMain.scala 28:24]
  wire [3:0] nutshell_io_frontend_awqos; // @[TopMain.scala 28:24]
  wire  nutshell_io_frontend_wready; // @[TopMain.scala 28:24]
  wire  nutshell_io_frontend_wvalid; // @[TopMain.scala 28:24]
  wire [63:0] nutshell_io_frontend_wdata; // @[TopMain.scala 28:24]
  wire [7:0] nutshell_io_frontend_wstrb; // @[TopMain.scala 28:24]
  wire  nutshell_io_frontend_wlast; // @[TopMain.scala 28:24]
  wire  nutshell_io_frontend_bready; // @[TopMain.scala 28:24]
  wire  nutshell_io_frontend_bvalid; // @[TopMain.scala 28:24]
  wire [1:0] nutshell_io_frontend_bresp; // @[TopMain.scala 28:24]
  wire  nutshell_io_frontend_bid; // @[TopMain.scala 28:24]
  wire  nutshell_io_frontend_buser; // @[TopMain.scala 28:24]
  wire  nutshell_io_frontend_arready; // @[TopMain.scala 28:24]
  wire  nutshell_io_frontend_arvalid; // @[TopMain.scala 28:24]
  wire [31:0] nutshell_io_frontend_araddr; // @[TopMain.scala 28:24]
  wire [2:0] nutshell_io_frontend_arprot; // @[TopMain.scala 28:24]
  wire  nutshell_io_frontend_arid; // @[TopMain.scala 28:24]
  wire  nutshell_io_frontend_aruser; // @[TopMain.scala 28:24]
  wire [7:0] nutshell_io_frontend_arlen; // @[TopMain.scala 28:24]
  wire [2:0] nutshell_io_frontend_arsize; // @[TopMain.scala 28:24]
  wire [1:0] nutshell_io_frontend_arburst; // @[TopMain.scala 28:24]
  wire  nutshell_io_frontend_arlock; // @[TopMain.scala 28:24]
  wire [3:0] nutshell_io_frontend_arcache; // @[TopMain.scala 28:24]
  wire [3:0] nutshell_io_frontend_arqos; // @[TopMain.scala 28:24]
  wire  nutshell_io_frontend_rready; // @[TopMain.scala 28:24]
  wire  nutshell_io_frontend_rvalid; // @[TopMain.scala 28:24]
  wire [1:0] nutshell_io_frontend_rresp; // @[TopMain.scala 28:24]
  wire [63:0] nutshell_io_frontend_rdata; // @[TopMain.scala 28:24]
  wire  nutshell_io_frontend_rlast; // @[TopMain.scala 28:24]
  wire  nutshell_io_frontend_rid; // @[TopMain.scala 28:24]
  wire  nutshell_io_frontend_ruser; // @[TopMain.scala 28:24]
  wire [2:0] nutshell_io_meip; // @[TopMain.scala 28:24]
  wire [38:0] nutshell_io_ila_WBUpc; // @[TopMain.scala 28:24]
  wire  nutshell_io_ila_WBUvalid; // @[TopMain.scala 28:24]
  wire  nutshell_io_ila_WBUrfWen; // @[TopMain.scala 28:24]
  wire [4:0] nutshell_io_ila_WBUrfDest; // @[TopMain.scala 28:24]
  wire [63:0] nutshell_io_ila_WBUrfData; // @[TopMain.scala 28:24]
  wire [63:0] nutshell_io_ila_InstrCnt; // @[TopMain.scala 28:24]
  wire  vga_clock; // @[TopMain.scala 29:19]
  wire  vga_reset; // @[TopMain.scala 29:19]
  wire  vga_io_in_fb_awready; // @[TopMain.scala 29:19]
  wire  vga_io_in_fb_awvalid; // @[TopMain.scala 29:19]
  wire [31:0] vga_io_in_fb_awaddr; // @[TopMain.scala 29:19]
  wire [2:0] vga_io_in_fb_awprot; // @[TopMain.scala 29:19]
  wire  vga_io_in_fb_wready; // @[TopMain.scala 29:19]
  wire  vga_io_in_fb_wvalid; // @[TopMain.scala 29:19]
  wire [63:0] vga_io_in_fb_wdata; // @[TopMain.scala 29:19]
  wire [7:0] vga_io_in_fb_wstrb; // @[TopMain.scala 29:19]
  wire  vga_io_in_fb_bready; // @[TopMain.scala 29:19]
  wire  vga_io_in_fb_bvalid; // @[TopMain.scala 29:19]
  wire [1:0] vga_io_in_fb_bresp; // @[TopMain.scala 29:19]
  wire  vga_io_in_fb_arready; // @[TopMain.scala 29:19]
  wire  vga_io_in_fb_arvalid; // @[TopMain.scala 29:19]
  wire [31:0] vga_io_in_fb_araddr; // @[TopMain.scala 29:19]
  wire [2:0] vga_io_in_fb_arprot; // @[TopMain.scala 29:19]
  wire  vga_io_in_fb_rready; // @[TopMain.scala 29:19]
  wire  vga_io_in_fb_rvalid; // @[TopMain.scala 29:19]
  wire [1:0] vga_io_in_fb_rresp; // @[TopMain.scala 29:19]
  wire [63:0] vga_io_in_fb_rdata; // @[TopMain.scala 29:19]
  wire  vga_io_in_ctrl_awready; // @[TopMain.scala 29:19]
  wire  vga_io_in_ctrl_awvalid; // @[TopMain.scala 29:19]
  wire [31:0] vga_io_in_ctrl_awaddr; // @[TopMain.scala 29:19]
  wire [2:0] vga_io_in_ctrl_awprot; // @[TopMain.scala 29:19]
  wire  vga_io_in_ctrl_wready; // @[TopMain.scala 29:19]
  wire  vga_io_in_ctrl_wvalid; // @[TopMain.scala 29:19]
  wire [63:0] vga_io_in_ctrl_wdata; // @[TopMain.scala 29:19]
  wire [7:0] vga_io_in_ctrl_wstrb; // @[TopMain.scala 29:19]
  wire  vga_io_in_ctrl_bready; // @[TopMain.scala 29:19]
  wire  vga_io_in_ctrl_bvalid; // @[TopMain.scala 29:19]
  wire [1:0] vga_io_in_ctrl_bresp; // @[TopMain.scala 29:19]
  wire  vga_io_in_ctrl_arready; // @[TopMain.scala 29:19]
  wire  vga_io_in_ctrl_arvalid; // @[TopMain.scala 29:19]
  wire [31:0] vga_io_in_ctrl_araddr; // @[TopMain.scala 29:19]
  wire [2:0] vga_io_in_ctrl_arprot; // @[TopMain.scala 29:19]
  wire  vga_io_in_ctrl_rready; // @[TopMain.scala 29:19]
  wire  vga_io_in_ctrl_rvalid; // @[TopMain.scala 29:19]
  wire [1:0] vga_io_in_ctrl_rresp; // @[TopMain.scala 29:19]
  wire [63:0] vga_io_in_ctrl_rdata; // @[TopMain.scala 29:19]
  wire [23:0] vga_io_vga_rgb; // @[TopMain.scala 29:19]
  wire  vga_io_vga_hsync; // @[TopMain.scala 29:19]
  wire  vga_io_vga_vsync; // @[TopMain.scala 29:19]
  wire  vga_io_vga_valid; // @[TopMain.scala 29:19]
  NutShell nutshell ( // @[TopMain.scala 28:24]
    .clock(nutshell_clock),
    .reset(nutshell_reset),
    .io_mem_awready(nutshell_io_mem_awready),
    .io_mem_awvalid(nutshell_io_mem_awvalid),
    .io_mem_awaddr(nutshell_io_mem_awaddr),
    .io_mem_awprot(nutshell_io_mem_awprot),
    .io_mem_awid(nutshell_io_mem_awid),
    .io_mem_awuser(nutshell_io_mem_awuser),
    .io_mem_awlen(nutshell_io_mem_awlen),
    .io_mem_awsize(nutshell_io_mem_awsize),
    .io_mem_awburst(nutshell_io_mem_awburst),
    .io_mem_awlock(nutshell_io_mem_awlock),
    .io_mem_awcache(nutshell_io_mem_awcache),
    .io_mem_awqos(nutshell_io_mem_awqos),
    .io_mem_wready(nutshell_io_mem_wready),
    .io_mem_wvalid(nutshell_io_mem_wvalid),
    .io_mem_wdata(nutshell_io_mem_wdata),
    .io_mem_wstrb(nutshell_io_mem_wstrb),
    .io_mem_wlast(nutshell_io_mem_wlast),
    .io_mem_bready(nutshell_io_mem_bready),
    .io_mem_bvalid(nutshell_io_mem_bvalid),
    .io_mem_bresp(nutshell_io_mem_bresp),
    .io_mem_bid(nutshell_io_mem_bid),
    .io_mem_buser(nutshell_io_mem_buser),
    .io_mem_arready(nutshell_io_mem_arready),
    .io_mem_arvalid(nutshell_io_mem_arvalid),
    .io_mem_araddr(nutshell_io_mem_araddr),
    .io_mem_arprot(nutshell_io_mem_arprot),
    .io_mem_arid(nutshell_io_mem_arid),
    .io_mem_aruser(nutshell_io_mem_aruser),
    .io_mem_arlen(nutshell_io_mem_arlen),
    .io_mem_arsize(nutshell_io_mem_arsize),
    .io_mem_arburst(nutshell_io_mem_arburst),
    .io_mem_arlock(nutshell_io_mem_arlock),
    .io_mem_arcache(nutshell_io_mem_arcache),
    .io_mem_arqos(nutshell_io_mem_arqos),
    .io_mem_rready(nutshell_io_mem_rready),
    .io_mem_rvalid(nutshell_io_mem_rvalid),
    .io_mem_rresp(nutshell_io_mem_rresp),
    .io_mem_rdata(nutshell_io_mem_rdata),
    .io_mem_rlast(nutshell_io_mem_rlast),
    .io_mem_rid(nutshell_io_mem_rid),
    .io_mem_ruser(nutshell_io_mem_ruser),
    .io_mmio_awready(nutshell_io_mmio_awready),
    .io_mmio_awvalid(nutshell_io_mmio_awvalid),
    .io_mmio_awaddr(nutshell_io_mmio_awaddr),
    .io_mmio_awprot(nutshell_io_mmio_awprot),
    .io_mmio_awid(nutshell_io_mmio_awid),
    .io_mmio_awuser(nutshell_io_mmio_awuser),
    .io_mmio_awlen(nutshell_io_mmio_awlen),
    .io_mmio_awsize(nutshell_io_mmio_awsize),
    .io_mmio_awburst(nutshell_io_mmio_awburst),
    .io_mmio_awlock(nutshell_io_mmio_awlock),
    .io_mmio_awcache(nutshell_io_mmio_awcache),
    .io_mmio_awqos(nutshell_io_mmio_awqos),
    .io_mmio_wready(nutshell_io_mmio_wready),
    .io_mmio_wvalid(nutshell_io_mmio_wvalid),
    .io_mmio_wdata(nutshell_io_mmio_wdata),
    .io_mmio_wstrb(nutshell_io_mmio_wstrb),
    .io_mmio_wlast(nutshell_io_mmio_wlast),
    .io_mmio_bready(nutshell_io_mmio_bready),
    .io_mmio_bvalid(nutshell_io_mmio_bvalid),
    .io_mmio_bresp(nutshell_io_mmio_bresp),
    .io_mmio_bid(nutshell_io_mmio_bid),
    .io_mmio_buser(nutshell_io_mmio_buser),
    .io_mmio_arready(nutshell_io_mmio_arready),
    .io_mmio_arvalid(nutshell_io_mmio_arvalid),
    .io_mmio_araddr(nutshell_io_mmio_araddr),
    .io_mmio_arprot(nutshell_io_mmio_arprot),
    .io_mmio_arid(nutshell_io_mmio_arid),
    .io_mmio_aruser(nutshell_io_mmio_aruser),
    .io_mmio_arlen(nutshell_io_mmio_arlen),
    .io_mmio_arsize(nutshell_io_mmio_arsize),
    .io_mmio_arburst(nutshell_io_mmio_arburst),
    .io_mmio_arlock(nutshell_io_mmio_arlock),
    .io_mmio_arcache(nutshell_io_mmio_arcache),
    .io_mmio_arqos(nutshell_io_mmio_arqos),
    .io_mmio_rready(nutshell_io_mmio_rready),
    .io_mmio_rvalid(nutshell_io_mmio_rvalid),
    .io_mmio_rresp(nutshell_io_mmio_rresp),
    .io_mmio_rdata(nutshell_io_mmio_rdata),
    .io_mmio_rlast(nutshell_io_mmio_rlast),
    .io_mmio_rid(nutshell_io_mmio_rid),
    .io_mmio_ruser(nutshell_io_mmio_ruser),
    .io_frontend_awready(nutshell_io_frontend_awready),
    .io_frontend_awvalid(nutshell_io_frontend_awvalid),
    .io_frontend_awaddr(nutshell_io_frontend_awaddr),
    .io_frontend_awprot(nutshell_io_frontend_awprot),
    .io_frontend_awid(nutshell_io_frontend_awid),
    .io_frontend_awuser(nutshell_io_frontend_awuser),
    .io_frontend_awlen(nutshell_io_frontend_awlen),
    .io_frontend_awsize(nutshell_io_frontend_awsize),
    .io_frontend_awburst(nutshell_io_frontend_awburst),
    .io_frontend_awlock(nutshell_io_frontend_awlock),
    .io_frontend_awcache(nutshell_io_frontend_awcache),
    .io_frontend_awqos(nutshell_io_frontend_awqos),
    .io_frontend_wready(nutshell_io_frontend_wready),
    .io_frontend_wvalid(nutshell_io_frontend_wvalid),
    .io_frontend_wdata(nutshell_io_frontend_wdata),
    .io_frontend_wstrb(nutshell_io_frontend_wstrb),
    .io_frontend_wlast(nutshell_io_frontend_wlast),
    .io_frontend_bready(nutshell_io_frontend_bready),
    .io_frontend_bvalid(nutshell_io_frontend_bvalid),
    .io_frontend_bresp(nutshell_io_frontend_bresp),
    .io_frontend_bid(nutshell_io_frontend_bid),
    .io_frontend_buser(nutshell_io_frontend_buser),
    .io_frontend_arready(nutshell_io_frontend_arready),
    .io_frontend_arvalid(nutshell_io_frontend_arvalid),
    .io_frontend_araddr(nutshell_io_frontend_araddr),
    .io_frontend_arprot(nutshell_io_frontend_arprot),
    .io_frontend_arid(nutshell_io_frontend_arid),
    .io_frontend_aruser(nutshell_io_frontend_aruser),
    .io_frontend_arlen(nutshell_io_frontend_arlen),
    .io_frontend_arsize(nutshell_io_frontend_arsize),
    .io_frontend_arburst(nutshell_io_frontend_arburst),
    .io_frontend_arlock(nutshell_io_frontend_arlock),
    .io_frontend_arcache(nutshell_io_frontend_arcache),
    .io_frontend_arqos(nutshell_io_frontend_arqos),
    .io_frontend_rready(nutshell_io_frontend_rready),
    .io_frontend_rvalid(nutshell_io_frontend_rvalid),
    .io_frontend_rresp(nutshell_io_frontend_rresp),
    .io_frontend_rdata(nutshell_io_frontend_rdata),
    .io_frontend_rlast(nutshell_io_frontend_rlast),
    .io_frontend_rid(nutshell_io_frontend_rid),
    .io_frontend_ruser(nutshell_io_frontend_ruser),
    .io_meip(nutshell_io_meip),
    .io_ila_WBUpc(nutshell_io_ila_WBUpc),
    .io_ila_WBUvalid(nutshell_io_ila_WBUvalid),
    .io_ila_WBUrfWen(nutshell_io_ila_WBUrfWen),
    .io_ila_WBUrfDest(nutshell_io_ila_WBUrfDest),
    .io_ila_WBUrfData(nutshell_io_ila_WBUrfData),
    .io_ila_InstrCnt(nutshell_io_ila_InstrCnt)
  );
  AXI4VGA vga ( // @[TopMain.scala 29:19]
    .clock(vga_clock),
    .reset(vga_reset),
    .io_in_fb_awready(vga_io_in_fb_awready),
    .io_in_fb_awvalid(vga_io_in_fb_awvalid),
    .io_in_fb_awaddr(vga_io_in_fb_awaddr),
    .io_in_fb_awprot(vga_io_in_fb_awprot),
    .io_in_fb_wready(vga_io_in_fb_wready),
    .io_in_fb_wvalid(vga_io_in_fb_wvalid),
    .io_in_fb_wdata(vga_io_in_fb_wdata),
    .io_in_fb_wstrb(vga_io_in_fb_wstrb),
    .io_in_fb_bready(vga_io_in_fb_bready),
    .io_in_fb_bvalid(vga_io_in_fb_bvalid),
    .io_in_fb_bresp(vga_io_in_fb_bresp),
    .io_in_fb_arready(vga_io_in_fb_arready),
    .io_in_fb_arvalid(vga_io_in_fb_arvalid),
    .io_in_fb_araddr(vga_io_in_fb_araddr),
    .io_in_fb_arprot(vga_io_in_fb_arprot),
    .io_in_fb_rready(vga_io_in_fb_rready),
    .io_in_fb_rvalid(vga_io_in_fb_rvalid),
    .io_in_fb_rresp(vga_io_in_fb_rresp),
    .io_in_fb_rdata(vga_io_in_fb_rdata),
    .io_in_ctrl_awready(vga_io_in_ctrl_awready),
    .io_in_ctrl_awvalid(vga_io_in_ctrl_awvalid),
    .io_in_ctrl_awaddr(vga_io_in_ctrl_awaddr),
    .io_in_ctrl_awprot(vga_io_in_ctrl_awprot),
    .io_in_ctrl_wready(vga_io_in_ctrl_wready),
    .io_in_ctrl_wvalid(vga_io_in_ctrl_wvalid),
    .io_in_ctrl_wdata(vga_io_in_ctrl_wdata),
    .io_in_ctrl_wstrb(vga_io_in_ctrl_wstrb),
    .io_in_ctrl_bready(vga_io_in_ctrl_bready),
    .io_in_ctrl_bvalid(vga_io_in_ctrl_bvalid),
    .io_in_ctrl_bresp(vga_io_in_ctrl_bresp),
    .io_in_ctrl_arready(vga_io_in_ctrl_arready),
    .io_in_ctrl_arvalid(vga_io_in_ctrl_arvalid),
    .io_in_ctrl_araddr(vga_io_in_ctrl_araddr),
    .io_in_ctrl_arprot(vga_io_in_ctrl_arprot),
    .io_in_ctrl_rready(vga_io_in_ctrl_rready),
    .io_in_ctrl_rvalid(vga_io_in_ctrl_rvalid),
    .io_in_ctrl_rresp(vga_io_in_ctrl_rresp),
    .io_in_ctrl_rdata(vga_io_in_ctrl_rdata),
    .io_vga_rgb(vga_io_vga_rgb),
    .io_vga_hsync(vga_io_vga_hsync),
    .io_vga_vsync(vga_io_vga_vsync),
    .io_vga_valid(vga_io_vga_valid)
  );
  assign nutshell_clock = clock;
  assign nutshell_reset = reset;
  assign nutshell_io_mem_awready = 1'h0;
  assign nutshell_io_mem_wready = 1'h0;
  assign nutshell_io_mem_bvalid = 1'h0;
  assign nutshell_io_mem_bresp = 2'h0;
  assign nutshell_io_mem_bid = 1'h0;
  assign nutshell_io_mem_buser = 1'h0;
  assign nutshell_io_mem_arready = 1'h0;
  assign nutshell_io_mem_rvalid = 1'h0;
  assign nutshell_io_mem_rresp = 2'h0;
  assign nutshell_io_mem_rdata = 64'h0;
  assign nutshell_io_mem_rlast = 1'h0;
  assign nutshell_io_mem_rid = 1'h0;
  assign nutshell_io_mem_ruser = 1'h0;
  assign nutshell_io_mmio_awready = 1'h0;
  assign nutshell_io_mmio_wready = 1'h0;
  assign nutshell_io_mmio_bvalid = 1'h0;
  assign nutshell_io_mmio_bresp = 2'h0;
  assign nutshell_io_mmio_bid = 1'h0;
  assign nutshell_io_mmio_buser = 1'h0;
  assign nutshell_io_mmio_arready = 1'h0;
  assign nutshell_io_mmio_rvalid = 1'h0;
  assign nutshell_io_mmio_rresp = 2'h0;
  assign nutshell_io_mmio_rdata = 64'h0;
  assign nutshell_io_mmio_rlast = 1'h0;
  assign nutshell_io_mmio_rid = 1'h0;
  assign nutshell_io_mmio_ruser = 1'h0;
  assign nutshell_io_frontend_awvalid = 1'h0;
  assign nutshell_io_frontend_awaddr = 32'h0;
  assign nutshell_io_frontend_awprot = 3'h0;
  assign nutshell_io_frontend_awid = 1'h0;
  assign nutshell_io_frontend_awuser = 1'h0;
  assign nutshell_io_frontend_awlen = 8'h0;
  assign nutshell_io_frontend_awsize = 3'h0;
  assign nutshell_io_frontend_awburst = 2'h0;
  assign nutshell_io_frontend_awlock = 1'h0;
  assign nutshell_io_frontend_awcache = 4'h0;
  assign nutshell_io_frontend_awqos = 4'h0;
  assign nutshell_io_frontend_wvalid = 1'h0;
  assign nutshell_io_frontend_wdata = 64'h0;
  assign nutshell_io_frontend_wstrb = 8'h0;
  assign nutshell_io_frontend_wlast = 1'h0;
  assign nutshell_io_frontend_bready = 1'h0;
  assign nutshell_io_frontend_arvalid = 1'h0;
  assign nutshell_io_frontend_araddr = 32'h0;
  assign nutshell_io_frontend_arprot = 3'h0;
  assign nutshell_io_frontend_arid = 1'h0;
  assign nutshell_io_frontend_aruser = 1'h0;
  assign nutshell_io_frontend_arlen = 8'h0;
  assign nutshell_io_frontend_arsize = 3'h0;
  assign nutshell_io_frontend_arburst = 2'h0;
  assign nutshell_io_frontend_arlock = 1'h0;
  assign nutshell_io_frontend_arcache = 4'h0;
  assign nutshell_io_frontend_arqos = 4'h0;
  assign nutshell_io_frontend_rready = 1'h0;
  assign nutshell_io_meip = 3'h0;
  assign vga_clock = clock;
  assign vga_reset = reset;
  assign vga_io_in_fb_awvalid = 1'h0;
  assign vga_io_in_fb_awaddr = 32'h0;
  assign vga_io_in_fb_awprot = 3'h0;
  assign vga_io_in_fb_wvalid = 1'h0;
  assign vga_io_in_fb_wdata = 64'h0;
  assign vga_io_in_fb_wstrb = 8'h0;
  assign vga_io_in_fb_bready = 1'h0;
  assign vga_io_in_fb_arvalid = 1'h0;
  assign vga_io_in_fb_araddr = 32'h0;
  assign vga_io_in_fb_arprot = 3'h0;
  assign vga_io_in_fb_rready = 1'h0;
  assign vga_io_in_ctrl_awvalid = 1'h0;
  assign vga_io_in_ctrl_awaddr = 32'h0;
  assign vga_io_in_ctrl_awprot = 3'h0;
  assign vga_io_in_ctrl_wvalid = 1'h0;
  assign vga_io_in_ctrl_wdata = 64'h0;
  assign vga_io_in_ctrl_wstrb = 8'h0;
  assign vga_io_in_ctrl_bready = 1'h0;
  assign vga_io_in_ctrl_arvalid = 1'h0;
  assign vga_io_in_ctrl_araddr = 32'h0;
  assign vga_io_in_ctrl_arprot = 3'h0;
  assign vga_io_in_ctrl_rready = 1'h0;
endmodule
module array(
  input  [8:0]  RW0_addr,
  input         RW0_en,
  input         RW0_clk,
  input         RW0_wmode,
  input  [72:0] RW0_wdata_0,
  output [72:0] RW0_rdata_0
);
  wire [8:0] array_ext_RW0_addr;
  wire  array_ext_RW0_en;
  wire  array_ext_RW0_clk;
  wire  array_ext_RW0_wmode;
  wire [72:0] array_ext_RW0_wdata;
  wire [72:0] array_ext_RW0_rdata;
  array_ext array_ext (
    .RW0_addr(array_ext_RW0_addr),
    .RW0_en(array_ext_RW0_en),
    .RW0_clk(array_ext_RW0_clk),
    .RW0_wmode(array_ext_RW0_wmode),
    .RW0_wdata(array_ext_RW0_wdata),
    .RW0_rdata(array_ext_RW0_rdata)
  );
  assign array_ext_RW0_clk = RW0_clk;
  assign array_ext_RW0_en = RW0_en;
  assign array_ext_RW0_addr = RW0_addr;
  assign RW0_rdata_0 = array_ext_RW0_rdata;
  assign array_ext_RW0_wmode = RW0_wmode;
  assign array_ext_RW0_wdata = RW0_wdata_0;
endmodule
module array_0(
  input  [6:0]  RW0_addr,
  input         RW0_en,
  input         RW0_clk,
  input         RW0_wmode,
  input  [20:0] RW0_wdata_0,
  input  [20:0] RW0_wdata_1,
  input  [20:0] RW0_wdata_2,
  input  [20:0] RW0_wdata_3,
  output [20:0] RW0_rdata_0,
  output [20:0] RW0_rdata_1,
  output [20:0] RW0_rdata_2,
  output [20:0] RW0_rdata_3,
  input         RW0_wmask_0,
  input         RW0_wmask_1,
  input         RW0_wmask_2,
  input         RW0_wmask_3
);
  wire [6:0] array_0_ext_RW0_addr;
  wire  array_0_ext_RW0_en;
  wire  array_0_ext_RW0_clk;
  wire  array_0_ext_RW0_wmode;
  wire [83:0] array_0_ext_RW0_wdata;
  wire [83:0] array_0_ext_RW0_rdata;
  wire [3:0] array_0_ext_RW0_wmask;
  wire [41:0] _GEN_0 = {RW0_wdata_3,RW0_wdata_2};
  wire [41:0] _GEN_1 = {RW0_wdata_1,RW0_wdata_0};
  wire [1:0] _GEN_2 = {RW0_wmask_3,RW0_wmask_2};
  wire [1:0] _GEN_3 = {RW0_wmask_1,RW0_wmask_0};
  array_0_ext array_0_ext (
    .RW0_addr(array_0_ext_RW0_addr),
    .RW0_en(array_0_ext_RW0_en),
    .RW0_clk(array_0_ext_RW0_clk),
    .RW0_wmode(array_0_ext_RW0_wmode),
    .RW0_wdata(array_0_ext_RW0_wdata),
    .RW0_rdata(array_0_ext_RW0_rdata),
    .RW0_wmask(array_0_ext_RW0_wmask)
  );
  assign array_0_ext_RW0_clk = RW0_clk;
  assign array_0_ext_RW0_en = RW0_en;
  assign array_0_ext_RW0_addr = RW0_addr;
  assign RW0_rdata_0 = array_0_ext_RW0_rdata[20:0];
  assign RW0_rdata_1 = array_0_ext_RW0_rdata[41:21];
  assign RW0_rdata_2 = array_0_ext_RW0_rdata[62:42];
  assign RW0_rdata_3 = array_0_ext_RW0_rdata[83:63];
  assign array_0_ext_RW0_wmode = RW0_wmode;
  assign array_0_ext_RW0_wdata = {_GEN_0,_GEN_1};
  assign array_0_ext_RW0_wmask = {_GEN_2,_GEN_3};
endmodule
module array_1(
  input  [9:0]  RW0_addr,
  input         RW0_en,
  input         RW0_clk,
  input         RW0_wmode,
  input  [63:0] RW0_wdata_0,
  input  [63:0] RW0_wdata_1,
  input  [63:0] RW0_wdata_2,
  input  [63:0] RW0_wdata_3,
  output [63:0] RW0_rdata_0,
  output [63:0] RW0_rdata_1,
  output [63:0] RW0_rdata_2,
  output [63:0] RW0_rdata_3,
  input         RW0_wmask_0,
  input         RW0_wmask_1,
  input         RW0_wmask_2,
  input         RW0_wmask_3
);
  wire [9:0] array_1_ext_RW0_addr;
  wire  array_1_ext_RW0_en;
  wire  array_1_ext_RW0_clk;
  wire  array_1_ext_RW0_wmode;
  wire [255:0] array_1_ext_RW0_wdata;
  wire [255:0] array_1_ext_RW0_rdata;
  wire [3:0] array_1_ext_RW0_wmask;
  wire [127:0] _GEN_0 = {RW0_wdata_3,RW0_wdata_2};
  wire [127:0] _GEN_1 = {RW0_wdata_1,RW0_wdata_0};
  wire [1:0] _GEN_2 = {RW0_wmask_3,RW0_wmask_2};
  wire [1:0] _GEN_3 = {RW0_wmask_1,RW0_wmask_0};
  array_1_ext array_1_ext (
    .RW0_addr(array_1_ext_RW0_addr),
    .RW0_en(array_1_ext_RW0_en),
    .RW0_clk(array_1_ext_RW0_clk),
    .RW0_wmode(array_1_ext_RW0_wmode),
    .RW0_wdata(array_1_ext_RW0_wdata),
    .RW0_rdata(array_1_ext_RW0_rdata),
    .RW0_wmask(array_1_ext_RW0_wmask)
  );
  assign array_1_ext_RW0_clk = RW0_clk;
  assign array_1_ext_RW0_en = RW0_en;
  assign array_1_ext_RW0_addr = RW0_addr;
  assign RW0_rdata_0 = array_1_ext_RW0_rdata[63:0];
  assign RW0_rdata_1 = array_1_ext_RW0_rdata[127:64];
  assign RW0_rdata_2 = array_1_ext_RW0_rdata[191:128];
  assign RW0_rdata_3 = array_1_ext_RW0_rdata[255:192];
  assign array_1_ext_RW0_wmode = RW0_wmode;
  assign array_1_ext_RW0_wdata = {_GEN_0,_GEN_1};
  assign array_1_ext_RW0_wmask = {_GEN_2,_GEN_3};
endmodule
module array_2(
  input  [8:0]  RW0_addr,
  input         RW0_en,
  input         RW0_clk,
  input         RW0_wmode,
  input  [18:0] RW0_wdata_0,
  input  [18:0] RW0_wdata_1,
  input  [18:0] RW0_wdata_2,
  input  [18:0] RW0_wdata_3,
  output [18:0] RW0_rdata_0,
  output [18:0] RW0_rdata_1,
  output [18:0] RW0_rdata_2,
  output [18:0] RW0_rdata_3,
  input         RW0_wmask_0,
  input         RW0_wmask_1,
  input         RW0_wmask_2,
  input         RW0_wmask_3
);
  wire [8:0] array_2_ext_RW0_addr;
  wire  array_2_ext_RW0_en;
  wire  array_2_ext_RW0_clk;
  wire  array_2_ext_RW0_wmode;
  wire [75:0] array_2_ext_RW0_wdata;
  wire [75:0] array_2_ext_RW0_rdata;
  wire [3:0] array_2_ext_RW0_wmask;
  wire [37:0] _GEN_0 = {RW0_wdata_3,RW0_wdata_2};
  wire [37:0] _GEN_1 = {RW0_wdata_1,RW0_wdata_0};
  wire [1:0] _GEN_2 = {RW0_wmask_3,RW0_wmask_2};
  wire [1:0] _GEN_3 = {RW0_wmask_1,RW0_wmask_0};
  array_2_ext array_2_ext (
    .RW0_addr(array_2_ext_RW0_addr),
    .RW0_en(array_2_ext_RW0_en),
    .RW0_clk(array_2_ext_RW0_clk),
    .RW0_wmode(array_2_ext_RW0_wmode),
    .RW0_wdata(array_2_ext_RW0_wdata),
    .RW0_rdata(array_2_ext_RW0_rdata),
    .RW0_wmask(array_2_ext_RW0_wmask)
  );
  assign array_2_ext_RW0_clk = RW0_clk;
  assign array_2_ext_RW0_en = RW0_en;
  assign array_2_ext_RW0_addr = RW0_addr;
  assign RW0_rdata_0 = array_2_ext_RW0_rdata[18:0];
  assign RW0_rdata_1 = array_2_ext_RW0_rdata[37:19];
  assign RW0_rdata_2 = array_2_ext_RW0_rdata[56:38];
  assign RW0_rdata_3 = array_2_ext_RW0_rdata[75:57];
  assign array_2_ext_RW0_wmode = RW0_wmode;
  assign array_2_ext_RW0_wdata = {_GEN_0,_GEN_1};
  assign array_2_ext_RW0_wmask = {_GEN_2,_GEN_3};
endmodule
module array_3(
  input  [11:0] RW0_addr,
  input         RW0_en,
  input         RW0_clk,
  input         RW0_wmode,
  input  [63:0] RW0_wdata_0,
  input  [63:0] RW0_wdata_1,
  input  [63:0] RW0_wdata_2,
  input  [63:0] RW0_wdata_3,
  output [63:0] RW0_rdata_0,
  output [63:0] RW0_rdata_1,
  output [63:0] RW0_rdata_2,
  output [63:0] RW0_rdata_3,
  input         RW0_wmask_0,
  input         RW0_wmask_1,
  input         RW0_wmask_2,
  input         RW0_wmask_3
);
  wire [11:0] array_3_ext_RW0_addr;
  wire  array_3_ext_RW0_en;
  wire  array_3_ext_RW0_clk;
  wire  array_3_ext_RW0_wmode;
  wire [255:0] array_3_ext_RW0_wdata;
  wire [255:0] array_3_ext_RW0_rdata;
  wire [3:0] array_3_ext_RW0_wmask;
  wire [127:0] _GEN_0 = {RW0_wdata_3,RW0_wdata_2};
  wire [127:0] _GEN_1 = {RW0_wdata_1,RW0_wdata_0};
  wire [1:0] _GEN_2 = {RW0_wmask_3,RW0_wmask_2};
  wire [1:0] _GEN_3 = {RW0_wmask_1,RW0_wmask_0};
  array_3_ext array_3_ext (
    .RW0_addr(array_3_ext_RW0_addr),
    .RW0_en(array_3_ext_RW0_en),
    .RW0_clk(array_3_ext_RW0_clk),
    .RW0_wmode(array_3_ext_RW0_wmode),
    .RW0_wdata(array_3_ext_RW0_wdata),
    .RW0_rdata(array_3_ext_RW0_rdata),
    .RW0_wmask(array_3_ext_RW0_wmask)
  );
  assign array_3_ext_RW0_clk = RW0_clk;
  assign array_3_ext_RW0_en = RW0_en;
  assign array_3_ext_RW0_addr = RW0_addr;
  assign RW0_rdata_0 = array_3_ext_RW0_rdata[63:0];
  assign RW0_rdata_1 = array_3_ext_RW0_rdata[127:64];
  assign RW0_rdata_2 = array_3_ext_RW0_rdata[191:128];
  assign RW0_rdata_3 = array_3_ext_RW0_rdata[255:192];
  assign array_3_ext_RW0_wmode = RW0_wmode;
  assign array_3_ext_RW0_wdata = {_GEN_0,_GEN_1};
  assign array_3_ext_RW0_wmask = {_GEN_2,_GEN_3};
endmodule

module array_ext(
  input RW0_clk,
  input [8:0] RW0_addr,
  input RW0_en,
  input RW0_wmode,
  input [72:0] RW0_wdata,
  output [72:0] RW0_rdata
);

  reg reg_RW0_ren;
  reg [8:0] reg_RW0_addr;
  reg [72:0] ram [511:0];
  `ifdef RANDOMIZE_MEM_INIT
    integer initvar;
    initial begin
      #`RANDOMIZE_DELAY begin end
      for (initvar = 0; initvar < 512; initvar = initvar+1)
        ram[initvar] = {3 {$random}};
      reg_RW0_addr = {1 {$random}};
    end
  `endif
  integer i;
  always @(posedge RW0_clk)
    reg_RW0_ren <= RW0_en && !RW0_wmode;
  always @(posedge RW0_clk)
    if (RW0_en && !RW0_wmode) reg_RW0_addr <= RW0_addr;
  always @(posedge RW0_clk)
    if (RW0_en && RW0_wmode) begin
      for(i=0;i<1;i=i+1) begin
        ram[RW0_addr][i*73 +: 73] <= RW0_wdata[i*73 +: 73];
      end
    end
  `ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [95:0] RW0_random;
  `ifdef RANDOMIZE_MEM_INIT
    initial begin
      #`RANDOMIZE_DELAY begin end
      RW0_random = {$random, $random, $random};
      reg_RW0_ren = RW0_random[0];
    end
  `endif
  always @(posedge RW0_clk) RW0_random <= {$random, $random, $random};
  assign RW0_rdata = reg_RW0_ren ? ram[reg_RW0_addr] : RW0_random[72:0];
  `else
  assign RW0_rdata = ram[reg_RW0_addr];
  `endif

endmodule

module array_0_ext(
  input RW0_clk,
  input [6:0] RW0_addr,
  input RW0_en,
  input RW0_wmode,
  input [3:0] RW0_wmask,
  input [83:0] RW0_wdata,
  output [83:0] RW0_rdata
);

  reg reg_RW0_ren;
  reg [6:0] reg_RW0_addr;
  reg [83:0] ram [127:0];
  `ifdef RANDOMIZE_MEM_INIT
    integer initvar;
    initial begin
      #`RANDOMIZE_DELAY begin end
      for (initvar = 0; initvar < 128; initvar = initvar+1)
        ram[initvar] = {3 {$random}};
      reg_RW0_addr = {1 {$random}};
    end
  `endif
  integer i;
  always @(posedge RW0_clk)
    reg_RW0_ren <= RW0_en && !RW0_wmode;
  always @(posedge RW0_clk)
    if (RW0_en && !RW0_wmode) reg_RW0_addr <= RW0_addr;
  always @(posedge RW0_clk)
    if (RW0_en && RW0_wmode) begin
      for(i=0;i<4;i=i+1) begin
        if(RW0_wmask[i]) begin
          ram[RW0_addr][i*21 +: 21] <= RW0_wdata[i*21 +: 21];
        end
      end
    end
  `ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [95:0] RW0_random;
  `ifdef RANDOMIZE_MEM_INIT
    initial begin
      #`RANDOMIZE_DELAY begin end
      RW0_random = {$random, $random, $random};
      reg_RW0_ren = RW0_random[0];
    end
  `endif
  always @(posedge RW0_clk) RW0_random <= {$random, $random, $random};
  assign RW0_rdata = reg_RW0_ren ? ram[reg_RW0_addr] : RW0_random[83:0];
  `else
  assign RW0_rdata = ram[reg_RW0_addr];
  `endif

endmodule

module array_1_ext(
  input RW0_clk,
  input [9:0] RW0_addr,
  input RW0_en,
  input RW0_wmode,
  input [3:0] RW0_wmask,
  input [255:0] RW0_wdata,
  output [255:0] RW0_rdata
);

  reg reg_RW0_ren;
  reg [9:0] reg_RW0_addr;
  reg [255:0] ram [1023:0];
  `ifdef RANDOMIZE_MEM_INIT
    integer initvar;
    initial begin
      #`RANDOMIZE_DELAY begin end
      for (initvar = 0; initvar < 1024; initvar = initvar+1)
        ram[initvar] = {8 {$random}};
      reg_RW0_addr = {1 {$random}};
    end
  `endif
  integer i;
  always @(posedge RW0_clk)
    reg_RW0_ren <= RW0_en && !RW0_wmode;
  always @(posedge RW0_clk)
    if (RW0_en && !RW0_wmode) reg_RW0_addr <= RW0_addr;
  always @(posedge RW0_clk)
    if (RW0_en && RW0_wmode) begin
      for(i=0;i<4;i=i+1) begin
        if(RW0_wmask[i]) begin
          ram[RW0_addr][i*64 +: 64] <= RW0_wdata[i*64 +: 64];
        end
      end
    end
  `ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [255:0] RW0_random;
  `ifdef RANDOMIZE_MEM_INIT
    initial begin
      #`RANDOMIZE_DELAY begin end
      RW0_random = {$random, $random, $random, $random, $random, $random, $random, $random};
      reg_RW0_ren = RW0_random[0];
    end
  `endif
  always @(posedge RW0_clk) RW0_random <= {$random, $random, $random, $random, $random, $random, $random, $random};
  assign RW0_rdata = reg_RW0_ren ? ram[reg_RW0_addr] : RW0_random[255:0];
  `else
  assign RW0_rdata = ram[reg_RW0_addr];
  `endif

endmodule

module array_2_ext(
  input RW0_clk,
  input [8:0] RW0_addr,
  input RW0_en,
  input RW0_wmode,
  input [3:0] RW0_wmask,
  input [75:0] RW0_wdata,
  output [75:0] RW0_rdata
);

  reg reg_RW0_ren;
  reg [8:0] reg_RW0_addr;
  reg [75:0] ram [511:0];
  `ifdef RANDOMIZE_MEM_INIT
    integer initvar;
    initial begin
      #`RANDOMIZE_DELAY begin end
      for (initvar = 0; initvar < 512; initvar = initvar+1)
        ram[initvar] = {3 {$random}};
      reg_RW0_addr = {1 {$random}};
    end
  `endif
  integer i;
  always @(posedge RW0_clk)
    reg_RW0_ren <= RW0_en && !RW0_wmode;
  always @(posedge RW0_clk)
    if (RW0_en && !RW0_wmode) reg_RW0_addr <= RW0_addr;
  always @(posedge RW0_clk)
    if (RW0_en && RW0_wmode) begin
      for(i=0;i<4;i=i+1) begin
        if(RW0_wmask[i]) begin
          ram[RW0_addr][i*19 +: 19] <= RW0_wdata[i*19 +: 19];
        end
      end
    end
  `ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [95:0] RW0_random;
  `ifdef RANDOMIZE_MEM_INIT
    initial begin
      #`RANDOMIZE_DELAY begin end
      RW0_random = {$random, $random, $random};
      reg_RW0_ren = RW0_random[0];
    end
  `endif
  always @(posedge RW0_clk) RW0_random <= {$random, $random, $random};
  assign RW0_rdata = reg_RW0_ren ? ram[reg_RW0_addr] : RW0_random[75:0];
  `else
  assign RW0_rdata = ram[reg_RW0_addr];
  `endif

endmodule

module array_3_ext(
  input RW0_clk,
  input [11:0] RW0_addr,
  input RW0_en,
  input RW0_wmode,
  input [3:0] RW0_wmask,
  input [255:0] RW0_wdata,
  output [255:0] RW0_rdata
);

  reg reg_RW0_ren;
  reg [11:0] reg_RW0_addr;
  reg [255:0] ram [4095:0];
  `ifdef RANDOMIZE_MEM_INIT
    integer initvar;
    initial begin
      #`RANDOMIZE_DELAY begin end
      for (initvar = 0; initvar < 4096; initvar = initvar+1)
        ram[initvar] = {8 {$random}};
      reg_RW0_addr = {1 {$random}};
    end
  `endif
  integer i;
  always @(posedge RW0_clk)
    reg_RW0_ren <= RW0_en && !RW0_wmode;
  always @(posedge RW0_clk)
    if (RW0_en && !RW0_wmode) reg_RW0_addr <= RW0_addr;
  always @(posedge RW0_clk)
    if (RW0_en && RW0_wmode) begin
      for(i=0;i<4;i=i+1) begin
        if(RW0_wmask[i]) begin
          ram[RW0_addr][i*64 +: 64] <= RW0_wdata[i*64 +: 64];
        end
      end
    end
  `ifdef RANDOMIZE_GARBAGE_ASSIGN
  reg [255:0] RW0_random;
  `ifdef RANDOMIZE_MEM_INIT
    initial begin
      #`RANDOMIZE_DELAY begin end
      RW0_random = {$random, $random, $random, $random, $random, $random, $random, $random};
      reg_RW0_ren = RW0_random[0];
    end
  `endif
  always @(posedge RW0_clk) RW0_random <= {$random, $random, $random, $random, $random, $random, $random, $random};
  assign RW0_rdata = reg_RW0_ren ? ram[reg_RW0_addr] : RW0_random[255:0];
  `else
  assign RW0_rdata = ram[reg_RW0_addr];
  `endif

endmodule
